`include "../src/booth_pkg.sv"
`include "../src/booth.sv"
`include "../src/dadda.sv"
`include "../src/fa.sv"
`include "../src/ha.sv"
`include "../src/multiplier.sv"
`include "../common/packet_in.sv"
`include "../common/packet_out.sv"
`include "../mbe/sequence_in.sv"
`include "../mbe/fsm_mbe.sv"
`include "../common/sequencer.sv"
`include "../common/driver.sv"
`include "../common/driver_out.sv"
`include "../common/monitor.sv"
`include "../common/monitor_out.sv"
`include "../common/agent.sv"
`include "../common/agent_out.sv"
`include "../mbe/refmod.sv"
`include "../common/comparator.sv"
`include "../common/env.sv"
`include "../common/simple_test.sv"
