/*--------------------------------------------------------------------------------*/
// Engineer: Simone Ruffini 	[simone.ruffini@studenti.polito.it],
//			 Marco Crisolgo 	[s305673@studenti.polito.it],
//			 Matteo Lago 		[s319914@studenti.polito.it],
//			 Renato Belmonte 	[s316792@studenti.polito.it],
//
// Module Name: Pipeline Register - DEC/EX
// Project Name: risc-v 
// Description: 
//
// Additional Comments: 
/*--------------------------------------------------------------------------------*/


module preg_dex_ex import riscv_pkg::*;
	(

    // control input signals
	input EX_ctrl EXctrl_in,
	input MEM_ctrl MEMctrl_in,
	input DEC_ctrl DECctrl_in, 

	// control output signals

    // data output signals

    // data input signals

);
    
endmodule
