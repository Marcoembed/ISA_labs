module fsm_mbe(dut_if.port_in in_inter, dut_if.port_out out_inter, output state_t state);

    always_ff @(posedge in_inter.clk)
    begin
        if(in_inter.rst) begin
            in_inter.ready <= 0;
            //out_inter.data <= 'x;
            out_inter.valid <= 0;
            state <= INITIAL;
        end
        else case(state)
                INITIAL: begin
                    in_inter.ready <= 1;
                    state <= WAIT;
                end
                
                WAIT: begin
                    if(in_inter.valid) begin
                        in_inter.ready <= 0;
                        //out_inter.data <= in_inter.A + in_inter.B;
                        $display("multiplier: input A = %d, input B = %d, output OUT = %d",in_inter.A[10:0],in_inter.B[10:0],out_inter.data);
                        $display("multiplier: input A = %b, input B = %b, output OUT = %b",in_inter.A[10:0],in_inter.B[10:0],out_inter.data);
                        out_inter.valid <= 1;
                        state <= SEND;
                    end
                end
                
                SEND: begin
                    if(out_inter.ready) begin
                        out_inter.valid <= 0;
                        in_inter.ready <= 1;
                        state <= WAIT;
                    end
                end
        endcase
    end
endmodule: fsm_mbe
