`include "../src/booth.sv"
`include "../src/dadda.sv"
`include "../src/fa.sv"
`include "../src/fpnew_classifier.sv"
`include "../src/fpnew_fma.sv"
`include "../src/fpnew_opgroup_block.sv"
`include "../src/fpnew_opgroup_fmt_slice.sv"
`include "../src/fpnew_rounding.sv"
`include "../src/fpnew_top.sv"
`include "../src/ha.sv"
`include "../src/lzc.sv"
`include "../src/multiplier.sv"
`include "../src/rr_arb_tree.sv"
`include "../common/packet_in.sv"
`include "../common/packet_out.sv"
`include "../fpm/sequence_in.sv"
`include "../fpm/fsm_fpm.sv"
`include "../common/sequencer.sv"
`include "../common/driver.sv"
`include "../common/driver_out.sv"
`include "../common/monitor.sv"
`include "../common/monitor_out.sv"
`include "../common/agent.sv"
`include "../common/agent_out.sv"
`include "../fpm/refmod.sv"
`include "../common/comparator.sv"
`include "../common/env.sv"
`include "../common/simple_test.sv"
