`include "../dadda/fa.sv"
`include "../dadda/ha.sv"

module dadda ();
	
// portmap

//ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

//ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

//ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

\\ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

\\ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

\\ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

\\ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

\\ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

\\ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

\\ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

\\ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

\\ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

\\ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

\\ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

\\ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

\\ITERATION: 0 Goal: 4

HA HA0_6 (pp[1][6], pp[2][4], s1[0][6], c1[0][7]);
HA HA0_7 (pp[1][7], pp[2][5], s1[0][7], c1[0][8]);
FA FA0_8 (pp[1][8], pp[2][6], pp[3][4], s1[0][8], c1[0][9]);
HA HA0_8 (pp[4][2], pp[5][0], s2[0][8], c2[0][9]);
FA FA0_9 (pp[1][9], pp[2][7], pp[3][5], s1[0][9], c1[0][10]);
HA HA0_9 (pp[4][3], pp[5][1], s2[0][9], c2[0][10]);
FA FA1_0_10 (pp[1][10], pp[2][8], pp[3][6], s1[0][10], c1[0][11]);
FA FA2_0_10 (pp[4][4], pp[5][2], pp[6][0], s2[0][10], c2[0][11]);
FA FA1_0_11 (b1, pp[2][9], pp[3][7], s1[0][11], c1[0][12]);
FA FA2_0_11 (pp[4][5], pp[5][3], pp[6][1], s2[0][11], c2[0][12]);
FA FA1_0_12 (b1, pp[2][10], pp[3][8], s1[0][12], c1[0][13]);
FA FA2_0_12 (pp[4][6], pp[5][4], pp[6][2], s2[0][12], c2[0][13]);
FA FA1_0_13 (!b1, !b3, pp[3][9], s1[0][13], c1[0][14]);
FA FA2_0_13 (pp[4][7], pp[5][5], pp[6][3], s2[0][13], c2[0][14]);
FA FA0_14 (1, pp[3][10], pp[4][8], s1[0][14], c1[0][15]);
HA HA0_14 (pp[5][6], pp[6][4], s2[0][14], c2[0][15]);
FA FA0_15 (!b5, pp[4][9], pp[5][7], s1[0][15], c1[0][16]);
HA HA0_16 (1, pp[4][10], s1[0][16], c1[0][17]);

\\ITERATION: 1 Goal: 3

HA HA1_4 (pp[1][4], pp[2][2], s1[1][4], c1[1][5]);
HA HA1_5 (pp[1][5], pp[2][3], s1[1][5], c1[1][6]);
FA FA1_6 (pp[3][2], pp[4][0], b7, s1[1][6], c1[1][7]);
FA FA1_7 (pp[3][3], pp[4][1], c1[0][7], s1[1][7], c1[1][8]);
FA FA1_8 (b9, c1[0][8], s1[0][8], s1[1][8], c1[1][9]);
FA FA1_9 (c1[0][9], c2[0][9], s1[0][9], s1[1][9], c1[1][10]);
FA FA1_10 (c1[0][10], c2[0][10], s1[0][10], s1[1][10], c1[1][11]);
FA FA1_11 (c1[0][11], c2[0][11], s1[0][11], s1[1][11], c1[1][12]);
FA FA1_12 (c1[0][12], c2[0][12], s1[0][12], s1[1][12], c1[1][13]);
FA FA1_13 (c1[0][13], c2[0][13], s1[0][13], s1[1][13], c1[1][14]);
FA FA1_14 (c1[0][14], c2[0][14], s1[0][14], s1[1][14], c1[1][15]);
FA FA1_15 (pp[6][5], c1[0][15], c2[0][15], s1[1][15], c1[1][16]);
FA FA1_16 (pp[5][8], pp[6][6], c1[0][16], s1[1][16], c1[1][17]);
FA FA1_17 (!b7, pp[5][9], pp[6][7], s1[1][17], c1[1][18]);
HA HA1_18 (1, pp[5][10], s1[1][18], c1[1][19]);

\\ITERATION: 2 Goal: 2

HA HA2_2 (pp[1][2], pp[2][0], s1[2][2], c1[2][3]);
HA HA2_3 (pp[1][3], pp[2][1], s1[2][3], c1[2][4]);
FA FA2_4 (pp[3][0], b5, s1[1][4], s1[2][4], c1[2][5]);
FA FA2_5 (pp[3][1], c1[1][5], s1[1][5], s1[2][5], c1[2][6]);
FA FA2_6 (s1[0][6], c1[1][6], s1[1][6], s1[2][6], c1[2][7]);
FA FA2_7 (s1[0][7], c1[1][7], s1[1][7], s1[2][7], c1[2][8]);
FA FA2_8 (s2[0][8], c1[1][8], s1[1][8], s1[2][8], c1[2][9]);
FA FA2_9 (s2[0][9], c1[1][9], s1[1][9], s1[2][9], c1[2][10]);
FA FA2_10 (s2[0][10], c1[1][10], s1[1][10], s1[2][10], c1[2][11]);
FA FA2_11 (s2[0][11], c1[1][11], s1[1][11], s1[2][11], c1[2][12]);
FA FA2_12 (s2[0][12], c1[1][12], s1[1][12], s1[2][12], c1[2][13]);
FA FA2_13 (s2[0][13], c1[1][13], s1[1][13], s1[2][13], c1[2][14]);
FA FA2_14 (s2[0][14], c1[1][14], s1[1][14], s1[2][14], c1[2][15]);
FA FA2_15 (s1[0][15], c1[1][15], s1[1][15], s1[2][15], c1[2][16]);
FA FA2_16 (s1[0][16], c1[1][16], s1[1][16], s1[2][16], c1[2][17]);
FA FA2_17 (c1[0][17], c1[1][17], s1[1][17], s1[2][17], c1[2][18]);
FA FA2_18 (pp[6][8], c1[1][18], s1[1][18], s1[2][18], c1[2][19]);
FA FA2_19 (!b9, pp[6][9], c1[1][19], s1[2][19], c1[2][20]);
// portmap

endmodule
