/*--------------------------------------------------------------------------------*/
// Engineer: Simone Ruffini 	[simone.ruffini@studenti.polito.it,
// 								 simoneruffini.work@gmail.com],
//			 Marco Crisolgo 	[s305673@studenti.polito.it],
//			 Matteo Lago 		[s319914@studenti.polito.it],
//			 Renato Belmonte 	[s316792@studenti.polito.it],
//
// Module Name: risc-v Datapath
// Project Name: risc-v 
// Description: 
//
// Additional Comments: 
/*--------------------------------------------------------------------------------*/

/*------------------------------*/
//	FETCH
/*------------------------------*/

/*------------------------------*/
//	DECODE
/*------------------------------*/

/*------------------------------*/
//	EXECUTE
/*------------------------------*/

/*------------------------------*/
//  MEMORY
/*------------------------------*/

/*------------------------------*/
//	WRITEBACK
/*------------------------------*/






