/*--------------------------------------------------------------------------------*/
// Engineer: Simone Ruffini 	[simone.ruffini@studenti.polito.it],
//			 Marco Crisolgo 	[s305673@studenti.polito.it],
//			 Matteo Lago 		[s319914@studenti.polito.it],
//			 Renato Belmonte 	[s316792@studenti.polito.it],
//
// Module Name: Control Unit
// Project Name: risc-v 
// Description: 
//
// Additional Comments: 
/*--------------------------------------------------------------------------------*/
import riscv_pkg::*;

module cu (
	input 	t_opcode opcode_i,
   	output 	EX_ctrl EX,	
   	output 	MEM_ctrl MEM,	
   	output 	WB_ctrl WB:	
);

always_comb begin 

end

endmodule


