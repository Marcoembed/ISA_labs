package dut_pkg;

typedef enum logic [1:0]{
    INITIAL,WAIT,SEND
} state_t;

endpackage: dut_pkg
