package booth_pkg;
		parameter pp_width 	= 11; 	//partial product number of bits
		parameter pp_deep	= 6;  	//number of partial prodcuts
		parameter level		= 2;  	//number of iteration levels
endpackage
	
