**************************************************
* OpenRAM generated memory.
* Words: 1024
* Data bits: 32
* Banks: 1
* Column mux: 8:1
**************************************************
* File: DFFPOSX1.pex.netlist
* Created: Wed Jan  2 18:36:24 2008
* Program "Calibre xRC"
* Version "v2007.2_34.24"
*
.subckt dff D Q clk vdd gnd
*
MM21 Q a_66_6# gnd gnd NMOS_VTG L=5e-08 W=5e-07
MM19 a_76_6# a_2_6# a_66_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM20 gnd Q a_76_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM18 a_66_6# clk a_61_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM17 a_61_6# a_34_4# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM10 gnd clk a_2_6# gnd NMOS_VTG L=5e-08 W=5e-07
MM16 a_34_4# a_22_6# gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM15 gnd a_34_4# a_31_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM14 a_31_6# clk a_22_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM13 a_22_6# a_2_6# a_17_6# gnd NMOS_VTG L=5e-08 W=2.5e-07
MM12 a_17_6# D gnd gnd NMOS_VTG L=5e-08 W=2.5e-07
MM11 Q a_66_6# vdd vdd PMOS_VTG L=5e-08 W=1e-06
MM9 vdd Q a_76_84# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM8 a_76_84# clk a_66_6# vdd PMOS_VTG L=5e-08 W=2.5e-07
MM7 a_66_6# a_2_6# a_61_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM6 a_61_74# a_34_4# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM0 vdd clk a_2_6# vdd PMOS_VTG L=5e-08 W=1e-06
MM5 a_34_4# a_22_6# vdd vdd PMOS_VTG L=5e-08 W=5e-07
MM4 vdd a_34_4# a_31_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM3 a_31_74# a_2_6# a_22_6# vdd PMOS_VTG L=5e-08 W=5e-07
MM2 a_22_6# clk a_17_74# vdd PMOS_VTG L=5e-08 W=5e-07
MM1 a_17_74# D vdd vdd PMOS_VTG L=5e-08 W=5e-07
* c_9 a_66_6# 0 0.271997f
* c_20 clk 0 0.350944f
* c_27 Q 0 0.202617f
* c_32 a_76_84# 0 0.0210573f
* c_38 a_76_6# 0 0.0204911f
* c_45 a_34_4# 0 0.172306f
* c_55 a_2_6# 0 0.283119f
* c_59 a_22_6# 0 0.157312f
* c_64 D 0 0.0816386f
* c_73 gnd 0 0.254131f
* c_81 vdd 0 0.23624f
*
*.include "dff.pex.netlist.dff.pxi"
*
.ends
*
*

.SUBCKT row_addr_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 7 cols: 1
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r1_c0 din_1 dout_1 clk vdd gnd dff
Xdff_r2_c0 din_2 dout_2 clk vdd gnd dff
Xdff_r3_c0 din_3 dout_3 clk vdd gnd dff
Xdff_r4_c0 din_4 dout_4 clk vdd gnd dff
Xdff_r5_c0 din_5 dout_5 clk vdd gnd dff
Xdff_r6_c0 din_6 dout_6 clk vdd gnd dff
.ENDS row_addr_dff

.SUBCKT col_addr_dff din_0 din_1 din_2 dout_0 dout_1 dout_2 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 3
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
.ENDS col_addr_dff

.SUBCKT data_dff din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 32
Xdff_r0_c0 din_0 dout_0 clk vdd gnd dff
Xdff_r0_c1 din_1 dout_1 clk vdd gnd dff
Xdff_r0_c2 din_2 dout_2 clk vdd gnd dff
Xdff_r0_c3 din_3 dout_3 clk vdd gnd dff
Xdff_r0_c4 din_4 dout_4 clk vdd gnd dff
Xdff_r0_c5 din_5 dout_5 clk vdd gnd dff
Xdff_r0_c6 din_6 dout_6 clk vdd gnd dff
Xdff_r0_c7 din_7 dout_7 clk vdd gnd dff
Xdff_r0_c8 din_8 dout_8 clk vdd gnd dff
Xdff_r0_c9 din_9 dout_9 clk vdd gnd dff
Xdff_r0_c10 din_10 dout_10 clk vdd gnd dff
Xdff_r0_c11 din_11 dout_11 clk vdd gnd dff
Xdff_r0_c12 din_12 dout_12 clk vdd gnd dff
Xdff_r0_c13 din_13 dout_13 clk vdd gnd dff
Xdff_r0_c14 din_14 dout_14 clk vdd gnd dff
Xdff_r0_c15 din_15 dout_15 clk vdd gnd dff
Xdff_r0_c16 din_16 dout_16 clk vdd gnd dff
Xdff_r0_c17 din_17 dout_17 clk vdd gnd dff
Xdff_r0_c18 din_18 dout_18 clk vdd gnd dff
Xdff_r0_c19 din_19 dout_19 clk vdd gnd dff
Xdff_r0_c20 din_20 dout_20 clk vdd gnd dff
Xdff_r0_c21 din_21 dout_21 clk vdd gnd dff
Xdff_r0_c22 din_22 dout_22 clk vdd gnd dff
Xdff_r0_c23 din_23 dout_23 clk vdd gnd dff
Xdff_r0_c24 din_24 dout_24 clk vdd gnd dff
Xdff_r0_c25 din_25 dout_25 clk vdd gnd dff
Xdff_r0_c26 din_26 dout_26 clk vdd gnd dff
Xdff_r0_c27 din_27 dout_27 clk vdd gnd dff
Xdff_r0_c28 din_28 dout_28 clk vdd gnd dff
Xdff_r0_c29 din_29 dout_29 clk vdd gnd dff
Xdff_r0_c30 din_30 dout_30 clk vdd gnd dff
Xdff_r0_c31 din_31 dout_31 clk vdd gnd dff
.ENDS data_dff

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT precharge_1 bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos1 bl en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mupper_pmos2 br en_bar vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS precharge_1

.SUBCKT precharge_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 bl_256 br_256 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* OUTPUT: bl_65 
* OUTPUT: br_65 
* OUTPUT: bl_66 
* OUTPUT: br_66 
* OUTPUT: bl_67 
* OUTPUT: br_67 
* OUTPUT: bl_68 
* OUTPUT: br_68 
* OUTPUT: bl_69 
* OUTPUT: br_69 
* OUTPUT: bl_70 
* OUTPUT: br_70 
* OUTPUT: bl_71 
* OUTPUT: br_71 
* OUTPUT: bl_72 
* OUTPUT: br_72 
* OUTPUT: bl_73 
* OUTPUT: br_73 
* OUTPUT: bl_74 
* OUTPUT: br_74 
* OUTPUT: bl_75 
* OUTPUT: br_75 
* OUTPUT: bl_76 
* OUTPUT: br_76 
* OUTPUT: bl_77 
* OUTPUT: br_77 
* OUTPUT: bl_78 
* OUTPUT: br_78 
* OUTPUT: bl_79 
* OUTPUT: br_79 
* OUTPUT: bl_80 
* OUTPUT: br_80 
* OUTPUT: bl_81 
* OUTPUT: br_81 
* OUTPUT: bl_82 
* OUTPUT: br_82 
* OUTPUT: bl_83 
* OUTPUT: br_83 
* OUTPUT: bl_84 
* OUTPUT: br_84 
* OUTPUT: bl_85 
* OUTPUT: br_85 
* OUTPUT: bl_86 
* OUTPUT: br_86 
* OUTPUT: bl_87 
* OUTPUT: br_87 
* OUTPUT: bl_88 
* OUTPUT: br_88 
* OUTPUT: bl_89 
* OUTPUT: br_89 
* OUTPUT: bl_90 
* OUTPUT: br_90 
* OUTPUT: bl_91 
* OUTPUT: br_91 
* OUTPUT: bl_92 
* OUTPUT: br_92 
* OUTPUT: bl_93 
* OUTPUT: br_93 
* OUTPUT: bl_94 
* OUTPUT: br_94 
* OUTPUT: bl_95 
* OUTPUT: br_95 
* OUTPUT: bl_96 
* OUTPUT: br_96 
* OUTPUT: bl_97 
* OUTPUT: br_97 
* OUTPUT: bl_98 
* OUTPUT: br_98 
* OUTPUT: bl_99 
* OUTPUT: br_99 
* OUTPUT: bl_100 
* OUTPUT: br_100 
* OUTPUT: bl_101 
* OUTPUT: br_101 
* OUTPUT: bl_102 
* OUTPUT: br_102 
* OUTPUT: bl_103 
* OUTPUT: br_103 
* OUTPUT: bl_104 
* OUTPUT: br_104 
* OUTPUT: bl_105 
* OUTPUT: br_105 
* OUTPUT: bl_106 
* OUTPUT: br_106 
* OUTPUT: bl_107 
* OUTPUT: br_107 
* OUTPUT: bl_108 
* OUTPUT: br_108 
* OUTPUT: bl_109 
* OUTPUT: br_109 
* OUTPUT: bl_110 
* OUTPUT: br_110 
* OUTPUT: bl_111 
* OUTPUT: br_111 
* OUTPUT: bl_112 
* OUTPUT: br_112 
* OUTPUT: bl_113 
* OUTPUT: br_113 
* OUTPUT: bl_114 
* OUTPUT: br_114 
* OUTPUT: bl_115 
* OUTPUT: br_115 
* OUTPUT: bl_116 
* OUTPUT: br_116 
* OUTPUT: bl_117 
* OUTPUT: br_117 
* OUTPUT: bl_118 
* OUTPUT: br_118 
* OUTPUT: bl_119 
* OUTPUT: br_119 
* OUTPUT: bl_120 
* OUTPUT: br_120 
* OUTPUT: bl_121 
* OUTPUT: br_121 
* OUTPUT: bl_122 
* OUTPUT: br_122 
* OUTPUT: bl_123 
* OUTPUT: br_123 
* OUTPUT: bl_124 
* OUTPUT: br_124 
* OUTPUT: bl_125 
* OUTPUT: br_125 
* OUTPUT: bl_126 
* OUTPUT: br_126 
* OUTPUT: bl_127 
* OUTPUT: br_127 
* OUTPUT: bl_128 
* OUTPUT: br_128 
* OUTPUT: bl_129 
* OUTPUT: br_129 
* OUTPUT: bl_130 
* OUTPUT: br_130 
* OUTPUT: bl_131 
* OUTPUT: br_131 
* OUTPUT: bl_132 
* OUTPUT: br_132 
* OUTPUT: bl_133 
* OUTPUT: br_133 
* OUTPUT: bl_134 
* OUTPUT: br_134 
* OUTPUT: bl_135 
* OUTPUT: br_135 
* OUTPUT: bl_136 
* OUTPUT: br_136 
* OUTPUT: bl_137 
* OUTPUT: br_137 
* OUTPUT: bl_138 
* OUTPUT: br_138 
* OUTPUT: bl_139 
* OUTPUT: br_139 
* OUTPUT: bl_140 
* OUTPUT: br_140 
* OUTPUT: bl_141 
* OUTPUT: br_141 
* OUTPUT: bl_142 
* OUTPUT: br_142 
* OUTPUT: bl_143 
* OUTPUT: br_143 
* OUTPUT: bl_144 
* OUTPUT: br_144 
* OUTPUT: bl_145 
* OUTPUT: br_145 
* OUTPUT: bl_146 
* OUTPUT: br_146 
* OUTPUT: bl_147 
* OUTPUT: br_147 
* OUTPUT: bl_148 
* OUTPUT: br_148 
* OUTPUT: bl_149 
* OUTPUT: br_149 
* OUTPUT: bl_150 
* OUTPUT: br_150 
* OUTPUT: bl_151 
* OUTPUT: br_151 
* OUTPUT: bl_152 
* OUTPUT: br_152 
* OUTPUT: bl_153 
* OUTPUT: br_153 
* OUTPUT: bl_154 
* OUTPUT: br_154 
* OUTPUT: bl_155 
* OUTPUT: br_155 
* OUTPUT: bl_156 
* OUTPUT: br_156 
* OUTPUT: bl_157 
* OUTPUT: br_157 
* OUTPUT: bl_158 
* OUTPUT: br_158 
* OUTPUT: bl_159 
* OUTPUT: br_159 
* OUTPUT: bl_160 
* OUTPUT: br_160 
* OUTPUT: bl_161 
* OUTPUT: br_161 
* OUTPUT: bl_162 
* OUTPUT: br_162 
* OUTPUT: bl_163 
* OUTPUT: br_163 
* OUTPUT: bl_164 
* OUTPUT: br_164 
* OUTPUT: bl_165 
* OUTPUT: br_165 
* OUTPUT: bl_166 
* OUTPUT: br_166 
* OUTPUT: bl_167 
* OUTPUT: br_167 
* OUTPUT: bl_168 
* OUTPUT: br_168 
* OUTPUT: bl_169 
* OUTPUT: br_169 
* OUTPUT: bl_170 
* OUTPUT: br_170 
* OUTPUT: bl_171 
* OUTPUT: br_171 
* OUTPUT: bl_172 
* OUTPUT: br_172 
* OUTPUT: bl_173 
* OUTPUT: br_173 
* OUTPUT: bl_174 
* OUTPUT: br_174 
* OUTPUT: bl_175 
* OUTPUT: br_175 
* OUTPUT: bl_176 
* OUTPUT: br_176 
* OUTPUT: bl_177 
* OUTPUT: br_177 
* OUTPUT: bl_178 
* OUTPUT: br_178 
* OUTPUT: bl_179 
* OUTPUT: br_179 
* OUTPUT: bl_180 
* OUTPUT: br_180 
* OUTPUT: bl_181 
* OUTPUT: br_181 
* OUTPUT: bl_182 
* OUTPUT: br_182 
* OUTPUT: bl_183 
* OUTPUT: br_183 
* OUTPUT: bl_184 
* OUTPUT: br_184 
* OUTPUT: bl_185 
* OUTPUT: br_185 
* OUTPUT: bl_186 
* OUTPUT: br_186 
* OUTPUT: bl_187 
* OUTPUT: br_187 
* OUTPUT: bl_188 
* OUTPUT: br_188 
* OUTPUT: bl_189 
* OUTPUT: br_189 
* OUTPUT: bl_190 
* OUTPUT: br_190 
* OUTPUT: bl_191 
* OUTPUT: br_191 
* OUTPUT: bl_192 
* OUTPUT: br_192 
* OUTPUT: bl_193 
* OUTPUT: br_193 
* OUTPUT: bl_194 
* OUTPUT: br_194 
* OUTPUT: bl_195 
* OUTPUT: br_195 
* OUTPUT: bl_196 
* OUTPUT: br_196 
* OUTPUT: bl_197 
* OUTPUT: br_197 
* OUTPUT: bl_198 
* OUTPUT: br_198 
* OUTPUT: bl_199 
* OUTPUT: br_199 
* OUTPUT: bl_200 
* OUTPUT: br_200 
* OUTPUT: bl_201 
* OUTPUT: br_201 
* OUTPUT: bl_202 
* OUTPUT: br_202 
* OUTPUT: bl_203 
* OUTPUT: br_203 
* OUTPUT: bl_204 
* OUTPUT: br_204 
* OUTPUT: bl_205 
* OUTPUT: br_205 
* OUTPUT: bl_206 
* OUTPUT: br_206 
* OUTPUT: bl_207 
* OUTPUT: br_207 
* OUTPUT: bl_208 
* OUTPUT: br_208 
* OUTPUT: bl_209 
* OUTPUT: br_209 
* OUTPUT: bl_210 
* OUTPUT: br_210 
* OUTPUT: bl_211 
* OUTPUT: br_211 
* OUTPUT: bl_212 
* OUTPUT: br_212 
* OUTPUT: bl_213 
* OUTPUT: br_213 
* OUTPUT: bl_214 
* OUTPUT: br_214 
* OUTPUT: bl_215 
* OUTPUT: br_215 
* OUTPUT: bl_216 
* OUTPUT: br_216 
* OUTPUT: bl_217 
* OUTPUT: br_217 
* OUTPUT: bl_218 
* OUTPUT: br_218 
* OUTPUT: bl_219 
* OUTPUT: br_219 
* OUTPUT: bl_220 
* OUTPUT: br_220 
* OUTPUT: bl_221 
* OUTPUT: br_221 
* OUTPUT: bl_222 
* OUTPUT: br_222 
* OUTPUT: bl_223 
* OUTPUT: br_223 
* OUTPUT: bl_224 
* OUTPUT: br_224 
* OUTPUT: bl_225 
* OUTPUT: br_225 
* OUTPUT: bl_226 
* OUTPUT: br_226 
* OUTPUT: bl_227 
* OUTPUT: br_227 
* OUTPUT: bl_228 
* OUTPUT: br_228 
* OUTPUT: bl_229 
* OUTPUT: br_229 
* OUTPUT: bl_230 
* OUTPUT: br_230 
* OUTPUT: bl_231 
* OUTPUT: br_231 
* OUTPUT: bl_232 
* OUTPUT: br_232 
* OUTPUT: bl_233 
* OUTPUT: br_233 
* OUTPUT: bl_234 
* OUTPUT: br_234 
* OUTPUT: bl_235 
* OUTPUT: br_235 
* OUTPUT: bl_236 
* OUTPUT: br_236 
* OUTPUT: bl_237 
* OUTPUT: br_237 
* OUTPUT: bl_238 
* OUTPUT: br_238 
* OUTPUT: bl_239 
* OUTPUT: br_239 
* OUTPUT: bl_240 
* OUTPUT: br_240 
* OUTPUT: bl_241 
* OUTPUT: br_241 
* OUTPUT: bl_242 
* OUTPUT: br_242 
* OUTPUT: bl_243 
* OUTPUT: br_243 
* OUTPUT: bl_244 
* OUTPUT: br_244 
* OUTPUT: bl_245 
* OUTPUT: br_245 
* OUTPUT: bl_246 
* OUTPUT: br_246 
* OUTPUT: bl_247 
* OUTPUT: br_247 
* OUTPUT: bl_248 
* OUTPUT: br_248 
* OUTPUT: bl_249 
* OUTPUT: br_249 
* OUTPUT: bl_250 
* OUTPUT: br_250 
* OUTPUT: bl_251 
* OUTPUT: br_251 
* OUTPUT: bl_252 
* OUTPUT: br_252 
* OUTPUT: bl_253 
* OUTPUT: br_253 
* OUTPUT: bl_254 
* OUTPUT: br_254 
* OUTPUT: bl_255 
* OUTPUT: br_255 
* OUTPUT: bl_256 
* OUTPUT: br_256 
* INPUT : en_bar 
* POWER : vdd 
* cols: 257 size: 1 bl: bl br: br
Xpre_column_0 bl_0 br_0 en_bar vdd precharge_1
Xpre_column_1 bl_1 br_1 en_bar vdd precharge_1
Xpre_column_2 bl_2 br_2 en_bar vdd precharge_1
Xpre_column_3 bl_3 br_3 en_bar vdd precharge_1
Xpre_column_4 bl_4 br_4 en_bar vdd precharge_1
Xpre_column_5 bl_5 br_5 en_bar vdd precharge_1
Xpre_column_6 bl_6 br_6 en_bar vdd precharge_1
Xpre_column_7 bl_7 br_7 en_bar vdd precharge_1
Xpre_column_8 bl_8 br_8 en_bar vdd precharge_1
Xpre_column_9 bl_9 br_9 en_bar vdd precharge_1
Xpre_column_10 bl_10 br_10 en_bar vdd precharge_1
Xpre_column_11 bl_11 br_11 en_bar vdd precharge_1
Xpre_column_12 bl_12 br_12 en_bar vdd precharge_1
Xpre_column_13 bl_13 br_13 en_bar vdd precharge_1
Xpre_column_14 bl_14 br_14 en_bar vdd precharge_1
Xpre_column_15 bl_15 br_15 en_bar vdd precharge_1
Xpre_column_16 bl_16 br_16 en_bar vdd precharge_1
Xpre_column_17 bl_17 br_17 en_bar vdd precharge_1
Xpre_column_18 bl_18 br_18 en_bar vdd precharge_1
Xpre_column_19 bl_19 br_19 en_bar vdd precharge_1
Xpre_column_20 bl_20 br_20 en_bar vdd precharge_1
Xpre_column_21 bl_21 br_21 en_bar vdd precharge_1
Xpre_column_22 bl_22 br_22 en_bar vdd precharge_1
Xpre_column_23 bl_23 br_23 en_bar vdd precharge_1
Xpre_column_24 bl_24 br_24 en_bar vdd precharge_1
Xpre_column_25 bl_25 br_25 en_bar vdd precharge_1
Xpre_column_26 bl_26 br_26 en_bar vdd precharge_1
Xpre_column_27 bl_27 br_27 en_bar vdd precharge_1
Xpre_column_28 bl_28 br_28 en_bar vdd precharge_1
Xpre_column_29 bl_29 br_29 en_bar vdd precharge_1
Xpre_column_30 bl_30 br_30 en_bar vdd precharge_1
Xpre_column_31 bl_31 br_31 en_bar vdd precharge_1
Xpre_column_32 bl_32 br_32 en_bar vdd precharge_1
Xpre_column_33 bl_33 br_33 en_bar vdd precharge_1
Xpre_column_34 bl_34 br_34 en_bar vdd precharge_1
Xpre_column_35 bl_35 br_35 en_bar vdd precharge_1
Xpre_column_36 bl_36 br_36 en_bar vdd precharge_1
Xpre_column_37 bl_37 br_37 en_bar vdd precharge_1
Xpre_column_38 bl_38 br_38 en_bar vdd precharge_1
Xpre_column_39 bl_39 br_39 en_bar vdd precharge_1
Xpre_column_40 bl_40 br_40 en_bar vdd precharge_1
Xpre_column_41 bl_41 br_41 en_bar vdd precharge_1
Xpre_column_42 bl_42 br_42 en_bar vdd precharge_1
Xpre_column_43 bl_43 br_43 en_bar vdd precharge_1
Xpre_column_44 bl_44 br_44 en_bar vdd precharge_1
Xpre_column_45 bl_45 br_45 en_bar vdd precharge_1
Xpre_column_46 bl_46 br_46 en_bar vdd precharge_1
Xpre_column_47 bl_47 br_47 en_bar vdd precharge_1
Xpre_column_48 bl_48 br_48 en_bar vdd precharge_1
Xpre_column_49 bl_49 br_49 en_bar vdd precharge_1
Xpre_column_50 bl_50 br_50 en_bar vdd precharge_1
Xpre_column_51 bl_51 br_51 en_bar vdd precharge_1
Xpre_column_52 bl_52 br_52 en_bar vdd precharge_1
Xpre_column_53 bl_53 br_53 en_bar vdd precharge_1
Xpre_column_54 bl_54 br_54 en_bar vdd precharge_1
Xpre_column_55 bl_55 br_55 en_bar vdd precharge_1
Xpre_column_56 bl_56 br_56 en_bar vdd precharge_1
Xpre_column_57 bl_57 br_57 en_bar vdd precharge_1
Xpre_column_58 bl_58 br_58 en_bar vdd precharge_1
Xpre_column_59 bl_59 br_59 en_bar vdd precharge_1
Xpre_column_60 bl_60 br_60 en_bar vdd precharge_1
Xpre_column_61 bl_61 br_61 en_bar vdd precharge_1
Xpre_column_62 bl_62 br_62 en_bar vdd precharge_1
Xpre_column_63 bl_63 br_63 en_bar vdd precharge_1
Xpre_column_64 bl_64 br_64 en_bar vdd precharge_1
Xpre_column_65 bl_65 br_65 en_bar vdd precharge_1
Xpre_column_66 bl_66 br_66 en_bar vdd precharge_1
Xpre_column_67 bl_67 br_67 en_bar vdd precharge_1
Xpre_column_68 bl_68 br_68 en_bar vdd precharge_1
Xpre_column_69 bl_69 br_69 en_bar vdd precharge_1
Xpre_column_70 bl_70 br_70 en_bar vdd precharge_1
Xpre_column_71 bl_71 br_71 en_bar vdd precharge_1
Xpre_column_72 bl_72 br_72 en_bar vdd precharge_1
Xpre_column_73 bl_73 br_73 en_bar vdd precharge_1
Xpre_column_74 bl_74 br_74 en_bar vdd precharge_1
Xpre_column_75 bl_75 br_75 en_bar vdd precharge_1
Xpre_column_76 bl_76 br_76 en_bar vdd precharge_1
Xpre_column_77 bl_77 br_77 en_bar vdd precharge_1
Xpre_column_78 bl_78 br_78 en_bar vdd precharge_1
Xpre_column_79 bl_79 br_79 en_bar vdd precharge_1
Xpre_column_80 bl_80 br_80 en_bar vdd precharge_1
Xpre_column_81 bl_81 br_81 en_bar vdd precharge_1
Xpre_column_82 bl_82 br_82 en_bar vdd precharge_1
Xpre_column_83 bl_83 br_83 en_bar vdd precharge_1
Xpre_column_84 bl_84 br_84 en_bar vdd precharge_1
Xpre_column_85 bl_85 br_85 en_bar vdd precharge_1
Xpre_column_86 bl_86 br_86 en_bar vdd precharge_1
Xpre_column_87 bl_87 br_87 en_bar vdd precharge_1
Xpre_column_88 bl_88 br_88 en_bar vdd precharge_1
Xpre_column_89 bl_89 br_89 en_bar vdd precharge_1
Xpre_column_90 bl_90 br_90 en_bar vdd precharge_1
Xpre_column_91 bl_91 br_91 en_bar vdd precharge_1
Xpre_column_92 bl_92 br_92 en_bar vdd precharge_1
Xpre_column_93 bl_93 br_93 en_bar vdd precharge_1
Xpre_column_94 bl_94 br_94 en_bar vdd precharge_1
Xpre_column_95 bl_95 br_95 en_bar vdd precharge_1
Xpre_column_96 bl_96 br_96 en_bar vdd precharge_1
Xpre_column_97 bl_97 br_97 en_bar vdd precharge_1
Xpre_column_98 bl_98 br_98 en_bar vdd precharge_1
Xpre_column_99 bl_99 br_99 en_bar vdd precharge_1
Xpre_column_100 bl_100 br_100 en_bar vdd precharge_1
Xpre_column_101 bl_101 br_101 en_bar vdd precharge_1
Xpre_column_102 bl_102 br_102 en_bar vdd precharge_1
Xpre_column_103 bl_103 br_103 en_bar vdd precharge_1
Xpre_column_104 bl_104 br_104 en_bar vdd precharge_1
Xpre_column_105 bl_105 br_105 en_bar vdd precharge_1
Xpre_column_106 bl_106 br_106 en_bar vdd precharge_1
Xpre_column_107 bl_107 br_107 en_bar vdd precharge_1
Xpre_column_108 bl_108 br_108 en_bar vdd precharge_1
Xpre_column_109 bl_109 br_109 en_bar vdd precharge_1
Xpre_column_110 bl_110 br_110 en_bar vdd precharge_1
Xpre_column_111 bl_111 br_111 en_bar vdd precharge_1
Xpre_column_112 bl_112 br_112 en_bar vdd precharge_1
Xpre_column_113 bl_113 br_113 en_bar vdd precharge_1
Xpre_column_114 bl_114 br_114 en_bar vdd precharge_1
Xpre_column_115 bl_115 br_115 en_bar vdd precharge_1
Xpre_column_116 bl_116 br_116 en_bar vdd precharge_1
Xpre_column_117 bl_117 br_117 en_bar vdd precharge_1
Xpre_column_118 bl_118 br_118 en_bar vdd precharge_1
Xpre_column_119 bl_119 br_119 en_bar vdd precharge_1
Xpre_column_120 bl_120 br_120 en_bar vdd precharge_1
Xpre_column_121 bl_121 br_121 en_bar vdd precharge_1
Xpre_column_122 bl_122 br_122 en_bar vdd precharge_1
Xpre_column_123 bl_123 br_123 en_bar vdd precharge_1
Xpre_column_124 bl_124 br_124 en_bar vdd precharge_1
Xpre_column_125 bl_125 br_125 en_bar vdd precharge_1
Xpre_column_126 bl_126 br_126 en_bar vdd precharge_1
Xpre_column_127 bl_127 br_127 en_bar vdd precharge_1
Xpre_column_128 bl_128 br_128 en_bar vdd precharge_1
Xpre_column_129 bl_129 br_129 en_bar vdd precharge_1
Xpre_column_130 bl_130 br_130 en_bar vdd precharge_1
Xpre_column_131 bl_131 br_131 en_bar vdd precharge_1
Xpre_column_132 bl_132 br_132 en_bar vdd precharge_1
Xpre_column_133 bl_133 br_133 en_bar vdd precharge_1
Xpre_column_134 bl_134 br_134 en_bar vdd precharge_1
Xpre_column_135 bl_135 br_135 en_bar vdd precharge_1
Xpre_column_136 bl_136 br_136 en_bar vdd precharge_1
Xpre_column_137 bl_137 br_137 en_bar vdd precharge_1
Xpre_column_138 bl_138 br_138 en_bar vdd precharge_1
Xpre_column_139 bl_139 br_139 en_bar vdd precharge_1
Xpre_column_140 bl_140 br_140 en_bar vdd precharge_1
Xpre_column_141 bl_141 br_141 en_bar vdd precharge_1
Xpre_column_142 bl_142 br_142 en_bar vdd precharge_1
Xpre_column_143 bl_143 br_143 en_bar vdd precharge_1
Xpre_column_144 bl_144 br_144 en_bar vdd precharge_1
Xpre_column_145 bl_145 br_145 en_bar vdd precharge_1
Xpre_column_146 bl_146 br_146 en_bar vdd precharge_1
Xpre_column_147 bl_147 br_147 en_bar vdd precharge_1
Xpre_column_148 bl_148 br_148 en_bar vdd precharge_1
Xpre_column_149 bl_149 br_149 en_bar vdd precharge_1
Xpre_column_150 bl_150 br_150 en_bar vdd precharge_1
Xpre_column_151 bl_151 br_151 en_bar vdd precharge_1
Xpre_column_152 bl_152 br_152 en_bar vdd precharge_1
Xpre_column_153 bl_153 br_153 en_bar vdd precharge_1
Xpre_column_154 bl_154 br_154 en_bar vdd precharge_1
Xpre_column_155 bl_155 br_155 en_bar vdd precharge_1
Xpre_column_156 bl_156 br_156 en_bar vdd precharge_1
Xpre_column_157 bl_157 br_157 en_bar vdd precharge_1
Xpre_column_158 bl_158 br_158 en_bar vdd precharge_1
Xpre_column_159 bl_159 br_159 en_bar vdd precharge_1
Xpre_column_160 bl_160 br_160 en_bar vdd precharge_1
Xpre_column_161 bl_161 br_161 en_bar vdd precharge_1
Xpre_column_162 bl_162 br_162 en_bar vdd precharge_1
Xpre_column_163 bl_163 br_163 en_bar vdd precharge_1
Xpre_column_164 bl_164 br_164 en_bar vdd precharge_1
Xpre_column_165 bl_165 br_165 en_bar vdd precharge_1
Xpre_column_166 bl_166 br_166 en_bar vdd precharge_1
Xpre_column_167 bl_167 br_167 en_bar vdd precharge_1
Xpre_column_168 bl_168 br_168 en_bar vdd precharge_1
Xpre_column_169 bl_169 br_169 en_bar vdd precharge_1
Xpre_column_170 bl_170 br_170 en_bar vdd precharge_1
Xpre_column_171 bl_171 br_171 en_bar vdd precharge_1
Xpre_column_172 bl_172 br_172 en_bar vdd precharge_1
Xpre_column_173 bl_173 br_173 en_bar vdd precharge_1
Xpre_column_174 bl_174 br_174 en_bar vdd precharge_1
Xpre_column_175 bl_175 br_175 en_bar vdd precharge_1
Xpre_column_176 bl_176 br_176 en_bar vdd precharge_1
Xpre_column_177 bl_177 br_177 en_bar vdd precharge_1
Xpre_column_178 bl_178 br_178 en_bar vdd precharge_1
Xpre_column_179 bl_179 br_179 en_bar vdd precharge_1
Xpre_column_180 bl_180 br_180 en_bar vdd precharge_1
Xpre_column_181 bl_181 br_181 en_bar vdd precharge_1
Xpre_column_182 bl_182 br_182 en_bar vdd precharge_1
Xpre_column_183 bl_183 br_183 en_bar vdd precharge_1
Xpre_column_184 bl_184 br_184 en_bar vdd precharge_1
Xpre_column_185 bl_185 br_185 en_bar vdd precharge_1
Xpre_column_186 bl_186 br_186 en_bar vdd precharge_1
Xpre_column_187 bl_187 br_187 en_bar vdd precharge_1
Xpre_column_188 bl_188 br_188 en_bar vdd precharge_1
Xpre_column_189 bl_189 br_189 en_bar vdd precharge_1
Xpre_column_190 bl_190 br_190 en_bar vdd precharge_1
Xpre_column_191 bl_191 br_191 en_bar vdd precharge_1
Xpre_column_192 bl_192 br_192 en_bar vdd precharge_1
Xpre_column_193 bl_193 br_193 en_bar vdd precharge_1
Xpre_column_194 bl_194 br_194 en_bar vdd precharge_1
Xpre_column_195 bl_195 br_195 en_bar vdd precharge_1
Xpre_column_196 bl_196 br_196 en_bar vdd precharge_1
Xpre_column_197 bl_197 br_197 en_bar vdd precharge_1
Xpre_column_198 bl_198 br_198 en_bar vdd precharge_1
Xpre_column_199 bl_199 br_199 en_bar vdd precharge_1
Xpre_column_200 bl_200 br_200 en_bar vdd precharge_1
Xpre_column_201 bl_201 br_201 en_bar vdd precharge_1
Xpre_column_202 bl_202 br_202 en_bar vdd precharge_1
Xpre_column_203 bl_203 br_203 en_bar vdd precharge_1
Xpre_column_204 bl_204 br_204 en_bar vdd precharge_1
Xpre_column_205 bl_205 br_205 en_bar vdd precharge_1
Xpre_column_206 bl_206 br_206 en_bar vdd precharge_1
Xpre_column_207 bl_207 br_207 en_bar vdd precharge_1
Xpre_column_208 bl_208 br_208 en_bar vdd precharge_1
Xpre_column_209 bl_209 br_209 en_bar vdd precharge_1
Xpre_column_210 bl_210 br_210 en_bar vdd precharge_1
Xpre_column_211 bl_211 br_211 en_bar vdd precharge_1
Xpre_column_212 bl_212 br_212 en_bar vdd precharge_1
Xpre_column_213 bl_213 br_213 en_bar vdd precharge_1
Xpre_column_214 bl_214 br_214 en_bar vdd precharge_1
Xpre_column_215 bl_215 br_215 en_bar vdd precharge_1
Xpre_column_216 bl_216 br_216 en_bar vdd precharge_1
Xpre_column_217 bl_217 br_217 en_bar vdd precharge_1
Xpre_column_218 bl_218 br_218 en_bar vdd precharge_1
Xpre_column_219 bl_219 br_219 en_bar vdd precharge_1
Xpre_column_220 bl_220 br_220 en_bar vdd precharge_1
Xpre_column_221 bl_221 br_221 en_bar vdd precharge_1
Xpre_column_222 bl_222 br_222 en_bar vdd precharge_1
Xpre_column_223 bl_223 br_223 en_bar vdd precharge_1
Xpre_column_224 bl_224 br_224 en_bar vdd precharge_1
Xpre_column_225 bl_225 br_225 en_bar vdd precharge_1
Xpre_column_226 bl_226 br_226 en_bar vdd precharge_1
Xpre_column_227 bl_227 br_227 en_bar vdd precharge_1
Xpre_column_228 bl_228 br_228 en_bar vdd precharge_1
Xpre_column_229 bl_229 br_229 en_bar vdd precharge_1
Xpre_column_230 bl_230 br_230 en_bar vdd precharge_1
Xpre_column_231 bl_231 br_231 en_bar vdd precharge_1
Xpre_column_232 bl_232 br_232 en_bar vdd precharge_1
Xpre_column_233 bl_233 br_233 en_bar vdd precharge_1
Xpre_column_234 bl_234 br_234 en_bar vdd precharge_1
Xpre_column_235 bl_235 br_235 en_bar vdd precharge_1
Xpre_column_236 bl_236 br_236 en_bar vdd precharge_1
Xpre_column_237 bl_237 br_237 en_bar vdd precharge_1
Xpre_column_238 bl_238 br_238 en_bar vdd precharge_1
Xpre_column_239 bl_239 br_239 en_bar vdd precharge_1
Xpre_column_240 bl_240 br_240 en_bar vdd precharge_1
Xpre_column_241 bl_241 br_241 en_bar vdd precharge_1
Xpre_column_242 bl_242 br_242 en_bar vdd precharge_1
Xpre_column_243 bl_243 br_243 en_bar vdd precharge_1
Xpre_column_244 bl_244 br_244 en_bar vdd precharge_1
Xpre_column_245 bl_245 br_245 en_bar vdd precharge_1
Xpre_column_246 bl_246 br_246 en_bar vdd precharge_1
Xpre_column_247 bl_247 br_247 en_bar vdd precharge_1
Xpre_column_248 bl_248 br_248 en_bar vdd precharge_1
Xpre_column_249 bl_249 br_249 en_bar vdd precharge_1
Xpre_column_250 bl_250 br_250 en_bar vdd precharge_1
Xpre_column_251 bl_251 br_251 en_bar vdd precharge_1
Xpre_column_252 bl_252 br_252 en_bar vdd precharge_1
Xpre_column_253 bl_253 br_253 en_bar vdd precharge_1
Xpre_column_254 bl_254 br_254 en_bar vdd precharge_1
Xpre_column_255 bl_255 br_255 en_bar vdd precharge_1
Xpre_column_256 bl_256 br_256 en_bar vdd precharge_1
.ENDS precharge_array_0

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sense_amp_array_0 data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3 data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 data_8 bl_8 br_8 data_9 bl_9 br_9 data_10 bl_10 br_10 data_11 bl_11 br_11 data_12 bl_12 br_12 data_13 bl_13 br_13 data_14 bl_14 br_14 data_15 bl_15 br_15 data_16 bl_16 br_16 data_17 bl_17 br_17 data_18 bl_18 br_18 data_19 bl_19 br_19 data_20 bl_20 br_20 data_21 bl_21 br_21 data_22 bl_22 br_22 data_23 bl_23 br_23 data_24 bl_24 br_24 data_25 bl_25 br_25 data_26 bl_26 br_26 data_27 bl_27 br_27 data_28 bl_28 br_28 data_29 bl_29 br_29 data_30 bl_30 br_30 data_31 bl_31 br_31 en vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* OUTPUT: data_8 
* INPUT : bl_8 
* INPUT : br_8 
* OUTPUT: data_9 
* INPUT : bl_9 
* INPUT : br_9 
* OUTPUT: data_10 
* INPUT : bl_10 
* INPUT : br_10 
* OUTPUT: data_11 
* INPUT : bl_11 
* INPUT : br_11 
* OUTPUT: data_12 
* INPUT : bl_12 
* INPUT : br_12 
* OUTPUT: data_13 
* INPUT : bl_13 
* INPUT : br_13 
* OUTPUT: data_14 
* INPUT : bl_14 
* INPUT : br_14 
* OUTPUT: data_15 
* INPUT : bl_15 
* INPUT : br_15 
* OUTPUT: data_16 
* INPUT : bl_16 
* INPUT : br_16 
* OUTPUT: data_17 
* INPUT : bl_17 
* INPUT : br_17 
* OUTPUT: data_18 
* INPUT : bl_18 
* INPUT : br_18 
* OUTPUT: data_19 
* INPUT : bl_19 
* INPUT : br_19 
* OUTPUT: data_20 
* INPUT : bl_20 
* INPUT : br_20 
* OUTPUT: data_21 
* INPUT : bl_21 
* INPUT : br_21 
* OUTPUT: data_22 
* INPUT : bl_22 
* INPUT : br_22 
* OUTPUT: data_23 
* INPUT : bl_23 
* INPUT : br_23 
* OUTPUT: data_24 
* INPUT : bl_24 
* INPUT : br_24 
* OUTPUT: data_25 
* INPUT : bl_25 
* INPUT : br_25 
* OUTPUT: data_26 
* INPUT : bl_26 
* INPUT : br_26 
* OUTPUT: data_27 
* INPUT : bl_27 
* INPUT : br_27 
* OUTPUT: data_28 
* INPUT : bl_28 
* INPUT : br_28 
* OUTPUT: data_29 
* INPUT : bl_29 
* INPUT : br_29 
* OUTPUT: data_30 
* INPUT : bl_30 
* INPUT : br_30 
* OUTPUT: data_31 
* INPUT : bl_31 
* INPUT : br_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* words_per_row: 8
Xsa_d0 bl_0 br_0 data_0 en vdd gnd sense_amp
Xsa_d1 bl_1 br_1 data_1 en vdd gnd sense_amp
Xsa_d2 bl_2 br_2 data_2 en vdd gnd sense_amp
Xsa_d3 bl_3 br_3 data_3 en vdd gnd sense_amp
Xsa_d4 bl_4 br_4 data_4 en vdd gnd sense_amp
Xsa_d5 bl_5 br_5 data_5 en vdd gnd sense_amp
Xsa_d6 bl_6 br_6 data_6 en vdd gnd sense_amp
Xsa_d7 bl_7 br_7 data_7 en vdd gnd sense_amp
Xsa_d8 bl_8 br_8 data_8 en vdd gnd sense_amp
Xsa_d9 bl_9 br_9 data_9 en vdd gnd sense_amp
Xsa_d10 bl_10 br_10 data_10 en vdd gnd sense_amp
Xsa_d11 bl_11 br_11 data_11 en vdd gnd sense_amp
Xsa_d12 bl_12 br_12 data_12 en vdd gnd sense_amp
Xsa_d13 bl_13 br_13 data_13 en vdd gnd sense_amp
Xsa_d14 bl_14 br_14 data_14 en vdd gnd sense_amp
Xsa_d15 bl_15 br_15 data_15 en vdd gnd sense_amp
Xsa_d16 bl_16 br_16 data_16 en vdd gnd sense_amp
Xsa_d17 bl_17 br_17 data_17 en vdd gnd sense_amp
Xsa_d18 bl_18 br_18 data_18 en vdd gnd sense_amp
Xsa_d19 bl_19 br_19 data_19 en vdd gnd sense_amp
Xsa_d20 bl_20 br_20 data_20 en vdd gnd sense_amp
Xsa_d21 bl_21 br_21 data_21 en vdd gnd sense_amp
Xsa_d22 bl_22 br_22 data_22 en vdd gnd sense_amp
Xsa_d23 bl_23 br_23 data_23 en vdd gnd sense_amp
Xsa_d24 bl_24 br_24 data_24 en vdd gnd sense_amp
Xsa_d25 bl_25 br_25 data_25 en vdd gnd sense_amp
Xsa_d26 bl_26 br_26 data_26 en vdd gnd sense_amp
Xsa_d27 bl_27 br_27 data_27 en vdd gnd sense_amp
Xsa_d28 bl_28 br_28 data_28 en vdd gnd sense_amp
Xsa_d29 bl_29 br_29 data_29 en vdd gnd sense_amp
Xsa_d30 bl_30 br_30 data_30 en vdd gnd sense_amp
Xsa_d31 bl_31 br_31 data_31 en vdd gnd sense_amp
.ENDS sense_amp_array_0

* ptx M{0} {1} nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT single_level_column_mux_0 bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Mmux_tx1 bl sel bl_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mmux_tx2 br sel br_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
.ENDS single_level_column_mux_0

.SUBCKT single_level_column_mux_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : sel_4 
* INOUT : sel_5 
* INOUT : sel_6 
* INOUT : sel_7 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : bl_out_8 
* INOUT : br_out_8 
* INOUT : bl_out_9 
* INOUT : br_out_9 
* INOUT : bl_out_10 
* INOUT : br_out_10 
* INOUT : bl_out_11 
* INOUT : br_out_11 
* INOUT : bl_out_12 
* INOUT : br_out_12 
* INOUT : bl_out_13 
* INOUT : br_out_13 
* INOUT : bl_out_14 
* INOUT : br_out_14 
* INOUT : bl_out_15 
* INOUT : br_out_15 
* INOUT : bl_out_16 
* INOUT : br_out_16 
* INOUT : bl_out_17 
* INOUT : br_out_17 
* INOUT : bl_out_18 
* INOUT : br_out_18 
* INOUT : bl_out_19 
* INOUT : br_out_19 
* INOUT : bl_out_20 
* INOUT : br_out_20 
* INOUT : bl_out_21 
* INOUT : br_out_21 
* INOUT : bl_out_22 
* INOUT : br_out_22 
* INOUT : bl_out_23 
* INOUT : br_out_23 
* INOUT : bl_out_24 
* INOUT : br_out_24 
* INOUT : bl_out_25 
* INOUT : br_out_25 
* INOUT : bl_out_26 
* INOUT : br_out_26 
* INOUT : bl_out_27 
* INOUT : br_out_27 
* INOUT : bl_out_28 
* INOUT : br_out_28 
* INOUT : bl_out_29 
* INOUT : br_out_29 
* INOUT : bl_out_30 
* INOUT : br_out_30 
* INOUT : bl_out_31 
* INOUT : br_out_31 
* INOUT : gnd 
* cols: 256 word_size: 32 bl: bl br: br
XXMUX0 bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd single_level_column_mux_0
XXMUX1 bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd single_level_column_mux_0
XXMUX2 bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd single_level_column_mux_0
XXMUX3 bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd single_level_column_mux_0
XXMUX4 bl_4 br_4 bl_out_0 br_out_0 sel_4 gnd single_level_column_mux_0
XXMUX5 bl_5 br_5 bl_out_0 br_out_0 sel_5 gnd single_level_column_mux_0
XXMUX6 bl_6 br_6 bl_out_0 br_out_0 sel_6 gnd single_level_column_mux_0
XXMUX7 bl_7 br_7 bl_out_0 br_out_0 sel_7 gnd single_level_column_mux_0
XXMUX8 bl_8 br_8 bl_out_1 br_out_1 sel_0 gnd single_level_column_mux_0
XXMUX9 bl_9 br_9 bl_out_1 br_out_1 sel_1 gnd single_level_column_mux_0
XXMUX10 bl_10 br_10 bl_out_1 br_out_1 sel_2 gnd single_level_column_mux_0
XXMUX11 bl_11 br_11 bl_out_1 br_out_1 sel_3 gnd single_level_column_mux_0
XXMUX12 bl_12 br_12 bl_out_1 br_out_1 sel_4 gnd single_level_column_mux_0
XXMUX13 bl_13 br_13 bl_out_1 br_out_1 sel_5 gnd single_level_column_mux_0
XXMUX14 bl_14 br_14 bl_out_1 br_out_1 sel_6 gnd single_level_column_mux_0
XXMUX15 bl_15 br_15 bl_out_1 br_out_1 sel_7 gnd single_level_column_mux_0
XXMUX16 bl_16 br_16 bl_out_2 br_out_2 sel_0 gnd single_level_column_mux_0
XXMUX17 bl_17 br_17 bl_out_2 br_out_2 sel_1 gnd single_level_column_mux_0
XXMUX18 bl_18 br_18 bl_out_2 br_out_2 sel_2 gnd single_level_column_mux_0
XXMUX19 bl_19 br_19 bl_out_2 br_out_2 sel_3 gnd single_level_column_mux_0
XXMUX20 bl_20 br_20 bl_out_2 br_out_2 sel_4 gnd single_level_column_mux_0
XXMUX21 bl_21 br_21 bl_out_2 br_out_2 sel_5 gnd single_level_column_mux_0
XXMUX22 bl_22 br_22 bl_out_2 br_out_2 sel_6 gnd single_level_column_mux_0
XXMUX23 bl_23 br_23 bl_out_2 br_out_2 sel_7 gnd single_level_column_mux_0
XXMUX24 bl_24 br_24 bl_out_3 br_out_3 sel_0 gnd single_level_column_mux_0
XXMUX25 bl_25 br_25 bl_out_3 br_out_3 sel_1 gnd single_level_column_mux_0
XXMUX26 bl_26 br_26 bl_out_3 br_out_3 sel_2 gnd single_level_column_mux_0
XXMUX27 bl_27 br_27 bl_out_3 br_out_3 sel_3 gnd single_level_column_mux_0
XXMUX28 bl_28 br_28 bl_out_3 br_out_3 sel_4 gnd single_level_column_mux_0
XXMUX29 bl_29 br_29 bl_out_3 br_out_3 sel_5 gnd single_level_column_mux_0
XXMUX30 bl_30 br_30 bl_out_3 br_out_3 sel_6 gnd single_level_column_mux_0
XXMUX31 bl_31 br_31 bl_out_3 br_out_3 sel_7 gnd single_level_column_mux_0
XXMUX32 bl_32 br_32 bl_out_4 br_out_4 sel_0 gnd single_level_column_mux_0
XXMUX33 bl_33 br_33 bl_out_4 br_out_4 sel_1 gnd single_level_column_mux_0
XXMUX34 bl_34 br_34 bl_out_4 br_out_4 sel_2 gnd single_level_column_mux_0
XXMUX35 bl_35 br_35 bl_out_4 br_out_4 sel_3 gnd single_level_column_mux_0
XXMUX36 bl_36 br_36 bl_out_4 br_out_4 sel_4 gnd single_level_column_mux_0
XXMUX37 bl_37 br_37 bl_out_4 br_out_4 sel_5 gnd single_level_column_mux_0
XXMUX38 bl_38 br_38 bl_out_4 br_out_4 sel_6 gnd single_level_column_mux_0
XXMUX39 bl_39 br_39 bl_out_4 br_out_4 sel_7 gnd single_level_column_mux_0
XXMUX40 bl_40 br_40 bl_out_5 br_out_5 sel_0 gnd single_level_column_mux_0
XXMUX41 bl_41 br_41 bl_out_5 br_out_5 sel_1 gnd single_level_column_mux_0
XXMUX42 bl_42 br_42 bl_out_5 br_out_5 sel_2 gnd single_level_column_mux_0
XXMUX43 bl_43 br_43 bl_out_5 br_out_5 sel_3 gnd single_level_column_mux_0
XXMUX44 bl_44 br_44 bl_out_5 br_out_5 sel_4 gnd single_level_column_mux_0
XXMUX45 bl_45 br_45 bl_out_5 br_out_5 sel_5 gnd single_level_column_mux_0
XXMUX46 bl_46 br_46 bl_out_5 br_out_5 sel_6 gnd single_level_column_mux_0
XXMUX47 bl_47 br_47 bl_out_5 br_out_5 sel_7 gnd single_level_column_mux_0
XXMUX48 bl_48 br_48 bl_out_6 br_out_6 sel_0 gnd single_level_column_mux_0
XXMUX49 bl_49 br_49 bl_out_6 br_out_6 sel_1 gnd single_level_column_mux_0
XXMUX50 bl_50 br_50 bl_out_6 br_out_6 sel_2 gnd single_level_column_mux_0
XXMUX51 bl_51 br_51 bl_out_6 br_out_6 sel_3 gnd single_level_column_mux_0
XXMUX52 bl_52 br_52 bl_out_6 br_out_6 sel_4 gnd single_level_column_mux_0
XXMUX53 bl_53 br_53 bl_out_6 br_out_6 sel_5 gnd single_level_column_mux_0
XXMUX54 bl_54 br_54 bl_out_6 br_out_6 sel_6 gnd single_level_column_mux_0
XXMUX55 bl_55 br_55 bl_out_6 br_out_6 sel_7 gnd single_level_column_mux_0
XXMUX56 bl_56 br_56 bl_out_7 br_out_7 sel_0 gnd single_level_column_mux_0
XXMUX57 bl_57 br_57 bl_out_7 br_out_7 sel_1 gnd single_level_column_mux_0
XXMUX58 bl_58 br_58 bl_out_7 br_out_7 sel_2 gnd single_level_column_mux_0
XXMUX59 bl_59 br_59 bl_out_7 br_out_7 sel_3 gnd single_level_column_mux_0
XXMUX60 bl_60 br_60 bl_out_7 br_out_7 sel_4 gnd single_level_column_mux_0
XXMUX61 bl_61 br_61 bl_out_7 br_out_7 sel_5 gnd single_level_column_mux_0
XXMUX62 bl_62 br_62 bl_out_7 br_out_7 sel_6 gnd single_level_column_mux_0
XXMUX63 bl_63 br_63 bl_out_7 br_out_7 sel_7 gnd single_level_column_mux_0
XXMUX64 bl_64 br_64 bl_out_8 br_out_8 sel_0 gnd single_level_column_mux_0
XXMUX65 bl_65 br_65 bl_out_8 br_out_8 sel_1 gnd single_level_column_mux_0
XXMUX66 bl_66 br_66 bl_out_8 br_out_8 sel_2 gnd single_level_column_mux_0
XXMUX67 bl_67 br_67 bl_out_8 br_out_8 sel_3 gnd single_level_column_mux_0
XXMUX68 bl_68 br_68 bl_out_8 br_out_8 sel_4 gnd single_level_column_mux_0
XXMUX69 bl_69 br_69 bl_out_8 br_out_8 sel_5 gnd single_level_column_mux_0
XXMUX70 bl_70 br_70 bl_out_8 br_out_8 sel_6 gnd single_level_column_mux_0
XXMUX71 bl_71 br_71 bl_out_8 br_out_8 sel_7 gnd single_level_column_mux_0
XXMUX72 bl_72 br_72 bl_out_9 br_out_9 sel_0 gnd single_level_column_mux_0
XXMUX73 bl_73 br_73 bl_out_9 br_out_9 sel_1 gnd single_level_column_mux_0
XXMUX74 bl_74 br_74 bl_out_9 br_out_9 sel_2 gnd single_level_column_mux_0
XXMUX75 bl_75 br_75 bl_out_9 br_out_9 sel_3 gnd single_level_column_mux_0
XXMUX76 bl_76 br_76 bl_out_9 br_out_9 sel_4 gnd single_level_column_mux_0
XXMUX77 bl_77 br_77 bl_out_9 br_out_9 sel_5 gnd single_level_column_mux_0
XXMUX78 bl_78 br_78 bl_out_9 br_out_9 sel_6 gnd single_level_column_mux_0
XXMUX79 bl_79 br_79 bl_out_9 br_out_9 sel_7 gnd single_level_column_mux_0
XXMUX80 bl_80 br_80 bl_out_10 br_out_10 sel_0 gnd single_level_column_mux_0
XXMUX81 bl_81 br_81 bl_out_10 br_out_10 sel_1 gnd single_level_column_mux_0
XXMUX82 bl_82 br_82 bl_out_10 br_out_10 sel_2 gnd single_level_column_mux_0
XXMUX83 bl_83 br_83 bl_out_10 br_out_10 sel_3 gnd single_level_column_mux_0
XXMUX84 bl_84 br_84 bl_out_10 br_out_10 sel_4 gnd single_level_column_mux_0
XXMUX85 bl_85 br_85 bl_out_10 br_out_10 sel_5 gnd single_level_column_mux_0
XXMUX86 bl_86 br_86 bl_out_10 br_out_10 sel_6 gnd single_level_column_mux_0
XXMUX87 bl_87 br_87 bl_out_10 br_out_10 sel_7 gnd single_level_column_mux_0
XXMUX88 bl_88 br_88 bl_out_11 br_out_11 sel_0 gnd single_level_column_mux_0
XXMUX89 bl_89 br_89 bl_out_11 br_out_11 sel_1 gnd single_level_column_mux_0
XXMUX90 bl_90 br_90 bl_out_11 br_out_11 sel_2 gnd single_level_column_mux_0
XXMUX91 bl_91 br_91 bl_out_11 br_out_11 sel_3 gnd single_level_column_mux_0
XXMUX92 bl_92 br_92 bl_out_11 br_out_11 sel_4 gnd single_level_column_mux_0
XXMUX93 bl_93 br_93 bl_out_11 br_out_11 sel_5 gnd single_level_column_mux_0
XXMUX94 bl_94 br_94 bl_out_11 br_out_11 sel_6 gnd single_level_column_mux_0
XXMUX95 bl_95 br_95 bl_out_11 br_out_11 sel_7 gnd single_level_column_mux_0
XXMUX96 bl_96 br_96 bl_out_12 br_out_12 sel_0 gnd single_level_column_mux_0
XXMUX97 bl_97 br_97 bl_out_12 br_out_12 sel_1 gnd single_level_column_mux_0
XXMUX98 bl_98 br_98 bl_out_12 br_out_12 sel_2 gnd single_level_column_mux_0
XXMUX99 bl_99 br_99 bl_out_12 br_out_12 sel_3 gnd single_level_column_mux_0
XXMUX100 bl_100 br_100 bl_out_12 br_out_12 sel_4 gnd single_level_column_mux_0
XXMUX101 bl_101 br_101 bl_out_12 br_out_12 sel_5 gnd single_level_column_mux_0
XXMUX102 bl_102 br_102 bl_out_12 br_out_12 sel_6 gnd single_level_column_mux_0
XXMUX103 bl_103 br_103 bl_out_12 br_out_12 sel_7 gnd single_level_column_mux_0
XXMUX104 bl_104 br_104 bl_out_13 br_out_13 sel_0 gnd single_level_column_mux_0
XXMUX105 bl_105 br_105 bl_out_13 br_out_13 sel_1 gnd single_level_column_mux_0
XXMUX106 bl_106 br_106 bl_out_13 br_out_13 sel_2 gnd single_level_column_mux_0
XXMUX107 bl_107 br_107 bl_out_13 br_out_13 sel_3 gnd single_level_column_mux_0
XXMUX108 bl_108 br_108 bl_out_13 br_out_13 sel_4 gnd single_level_column_mux_0
XXMUX109 bl_109 br_109 bl_out_13 br_out_13 sel_5 gnd single_level_column_mux_0
XXMUX110 bl_110 br_110 bl_out_13 br_out_13 sel_6 gnd single_level_column_mux_0
XXMUX111 bl_111 br_111 bl_out_13 br_out_13 sel_7 gnd single_level_column_mux_0
XXMUX112 bl_112 br_112 bl_out_14 br_out_14 sel_0 gnd single_level_column_mux_0
XXMUX113 bl_113 br_113 bl_out_14 br_out_14 sel_1 gnd single_level_column_mux_0
XXMUX114 bl_114 br_114 bl_out_14 br_out_14 sel_2 gnd single_level_column_mux_0
XXMUX115 bl_115 br_115 bl_out_14 br_out_14 sel_3 gnd single_level_column_mux_0
XXMUX116 bl_116 br_116 bl_out_14 br_out_14 sel_4 gnd single_level_column_mux_0
XXMUX117 bl_117 br_117 bl_out_14 br_out_14 sel_5 gnd single_level_column_mux_0
XXMUX118 bl_118 br_118 bl_out_14 br_out_14 sel_6 gnd single_level_column_mux_0
XXMUX119 bl_119 br_119 bl_out_14 br_out_14 sel_7 gnd single_level_column_mux_0
XXMUX120 bl_120 br_120 bl_out_15 br_out_15 sel_0 gnd single_level_column_mux_0
XXMUX121 bl_121 br_121 bl_out_15 br_out_15 sel_1 gnd single_level_column_mux_0
XXMUX122 bl_122 br_122 bl_out_15 br_out_15 sel_2 gnd single_level_column_mux_0
XXMUX123 bl_123 br_123 bl_out_15 br_out_15 sel_3 gnd single_level_column_mux_0
XXMUX124 bl_124 br_124 bl_out_15 br_out_15 sel_4 gnd single_level_column_mux_0
XXMUX125 bl_125 br_125 bl_out_15 br_out_15 sel_5 gnd single_level_column_mux_0
XXMUX126 bl_126 br_126 bl_out_15 br_out_15 sel_6 gnd single_level_column_mux_0
XXMUX127 bl_127 br_127 bl_out_15 br_out_15 sel_7 gnd single_level_column_mux_0
XXMUX128 bl_128 br_128 bl_out_16 br_out_16 sel_0 gnd single_level_column_mux_0
XXMUX129 bl_129 br_129 bl_out_16 br_out_16 sel_1 gnd single_level_column_mux_0
XXMUX130 bl_130 br_130 bl_out_16 br_out_16 sel_2 gnd single_level_column_mux_0
XXMUX131 bl_131 br_131 bl_out_16 br_out_16 sel_3 gnd single_level_column_mux_0
XXMUX132 bl_132 br_132 bl_out_16 br_out_16 sel_4 gnd single_level_column_mux_0
XXMUX133 bl_133 br_133 bl_out_16 br_out_16 sel_5 gnd single_level_column_mux_0
XXMUX134 bl_134 br_134 bl_out_16 br_out_16 sel_6 gnd single_level_column_mux_0
XXMUX135 bl_135 br_135 bl_out_16 br_out_16 sel_7 gnd single_level_column_mux_0
XXMUX136 bl_136 br_136 bl_out_17 br_out_17 sel_0 gnd single_level_column_mux_0
XXMUX137 bl_137 br_137 bl_out_17 br_out_17 sel_1 gnd single_level_column_mux_0
XXMUX138 bl_138 br_138 bl_out_17 br_out_17 sel_2 gnd single_level_column_mux_0
XXMUX139 bl_139 br_139 bl_out_17 br_out_17 sel_3 gnd single_level_column_mux_0
XXMUX140 bl_140 br_140 bl_out_17 br_out_17 sel_4 gnd single_level_column_mux_0
XXMUX141 bl_141 br_141 bl_out_17 br_out_17 sel_5 gnd single_level_column_mux_0
XXMUX142 bl_142 br_142 bl_out_17 br_out_17 sel_6 gnd single_level_column_mux_0
XXMUX143 bl_143 br_143 bl_out_17 br_out_17 sel_7 gnd single_level_column_mux_0
XXMUX144 bl_144 br_144 bl_out_18 br_out_18 sel_0 gnd single_level_column_mux_0
XXMUX145 bl_145 br_145 bl_out_18 br_out_18 sel_1 gnd single_level_column_mux_0
XXMUX146 bl_146 br_146 bl_out_18 br_out_18 sel_2 gnd single_level_column_mux_0
XXMUX147 bl_147 br_147 bl_out_18 br_out_18 sel_3 gnd single_level_column_mux_0
XXMUX148 bl_148 br_148 bl_out_18 br_out_18 sel_4 gnd single_level_column_mux_0
XXMUX149 bl_149 br_149 bl_out_18 br_out_18 sel_5 gnd single_level_column_mux_0
XXMUX150 bl_150 br_150 bl_out_18 br_out_18 sel_6 gnd single_level_column_mux_0
XXMUX151 bl_151 br_151 bl_out_18 br_out_18 sel_7 gnd single_level_column_mux_0
XXMUX152 bl_152 br_152 bl_out_19 br_out_19 sel_0 gnd single_level_column_mux_0
XXMUX153 bl_153 br_153 bl_out_19 br_out_19 sel_1 gnd single_level_column_mux_0
XXMUX154 bl_154 br_154 bl_out_19 br_out_19 sel_2 gnd single_level_column_mux_0
XXMUX155 bl_155 br_155 bl_out_19 br_out_19 sel_3 gnd single_level_column_mux_0
XXMUX156 bl_156 br_156 bl_out_19 br_out_19 sel_4 gnd single_level_column_mux_0
XXMUX157 bl_157 br_157 bl_out_19 br_out_19 sel_5 gnd single_level_column_mux_0
XXMUX158 bl_158 br_158 bl_out_19 br_out_19 sel_6 gnd single_level_column_mux_0
XXMUX159 bl_159 br_159 bl_out_19 br_out_19 sel_7 gnd single_level_column_mux_0
XXMUX160 bl_160 br_160 bl_out_20 br_out_20 sel_0 gnd single_level_column_mux_0
XXMUX161 bl_161 br_161 bl_out_20 br_out_20 sel_1 gnd single_level_column_mux_0
XXMUX162 bl_162 br_162 bl_out_20 br_out_20 sel_2 gnd single_level_column_mux_0
XXMUX163 bl_163 br_163 bl_out_20 br_out_20 sel_3 gnd single_level_column_mux_0
XXMUX164 bl_164 br_164 bl_out_20 br_out_20 sel_4 gnd single_level_column_mux_0
XXMUX165 bl_165 br_165 bl_out_20 br_out_20 sel_5 gnd single_level_column_mux_0
XXMUX166 bl_166 br_166 bl_out_20 br_out_20 sel_6 gnd single_level_column_mux_0
XXMUX167 bl_167 br_167 bl_out_20 br_out_20 sel_7 gnd single_level_column_mux_0
XXMUX168 bl_168 br_168 bl_out_21 br_out_21 sel_0 gnd single_level_column_mux_0
XXMUX169 bl_169 br_169 bl_out_21 br_out_21 sel_1 gnd single_level_column_mux_0
XXMUX170 bl_170 br_170 bl_out_21 br_out_21 sel_2 gnd single_level_column_mux_0
XXMUX171 bl_171 br_171 bl_out_21 br_out_21 sel_3 gnd single_level_column_mux_0
XXMUX172 bl_172 br_172 bl_out_21 br_out_21 sel_4 gnd single_level_column_mux_0
XXMUX173 bl_173 br_173 bl_out_21 br_out_21 sel_5 gnd single_level_column_mux_0
XXMUX174 bl_174 br_174 bl_out_21 br_out_21 sel_6 gnd single_level_column_mux_0
XXMUX175 bl_175 br_175 bl_out_21 br_out_21 sel_7 gnd single_level_column_mux_0
XXMUX176 bl_176 br_176 bl_out_22 br_out_22 sel_0 gnd single_level_column_mux_0
XXMUX177 bl_177 br_177 bl_out_22 br_out_22 sel_1 gnd single_level_column_mux_0
XXMUX178 bl_178 br_178 bl_out_22 br_out_22 sel_2 gnd single_level_column_mux_0
XXMUX179 bl_179 br_179 bl_out_22 br_out_22 sel_3 gnd single_level_column_mux_0
XXMUX180 bl_180 br_180 bl_out_22 br_out_22 sel_4 gnd single_level_column_mux_0
XXMUX181 bl_181 br_181 bl_out_22 br_out_22 sel_5 gnd single_level_column_mux_0
XXMUX182 bl_182 br_182 bl_out_22 br_out_22 sel_6 gnd single_level_column_mux_0
XXMUX183 bl_183 br_183 bl_out_22 br_out_22 sel_7 gnd single_level_column_mux_0
XXMUX184 bl_184 br_184 bl_out_23 br_out_23 sel_0 gnd single_level_column_mux_0
XXMUX185 bl_185 br_185 bl_out_23 br_out_23 sel_1 gnd single_level_column_mux_0
XXMUX186 bl_186 br_186 bl_out_23 br_out_23 sel_2 gnd single_level_column_mux_0
XXMUX187 bl_187 br_187 bl_out_23 br_out_23 sel_3 gnd single_level_column_mux_0
XXMUX188 bl_188 br_188 bl_out_23 br_out_23 sel_4 gnd single_level_column_mux_0
XXMUX189 bl_189 br_189 bl_out_23 br_out_23 sel_5 gnd single_level_column_mux_0
XXMUX190 bl_190 br_190 bl_out_23 br_out_23 sel_6 gnd single_level_column_mux_0
XXMUX191 bl_191 br_191 bl_out_23 br_out_23 sel_7 gnd single_level_column_mux_0
XXMUX192 bl_192 br_192 bl_out_24 br_out_24 sel_0 gnd single_level_column_mux_0
XXMUX193 bl_193 br_193 bl_out_24 br_out_24 sel_1 gnd single_level_column_mux_0
XXMUX194 bl_194 br_194 bl_out_24 br_out_24 sel_2 gnd single_level_column_mux_0
XXMUX195 bl_195 br_195 bl_out_24 br_out_24 sel_3 gnd single_level_column_mux_0
XXMUX196 bl_196 br_196 bl_out_24 br_out_24 sel_4 gnd single_level_column_mux_0
XXMUX197 bl_197 br_197 bl_out_24 br_out_24 sel_5 gnd single_level_column_mux_0
XXMUX198 bl_198 br_198 bl_out_24 br_out_24 sel_6 gnd single_level_column_mux_0
XXMUX199 bl_199 br_199 bl_out_24 br_out_24 sel_7 gnd single_level_column_mux_0
XXMUX200 bl_200 br_200 bl_out_25 br_out_25 sel_0 gnd single_level_column_mux_0
XXMUX201 bl_201 br_201 bl_out_25 br_out_25 sel_1 gnd single_level_column_mux_0
XXMUX202 bl_202 br_202 bl_out_25 br_out_25 sel_2 gnd single_level_column_mux_0
XXMUX203 bl_203 br_203 bl_out_25 br_out_25 sel_3 gnd single_level_column_mux_0
XXMUX204 bl_204 br_204 bl_out_25 br_out_25 sel_4 gnd single_level_column_mux_0
XXMUX205 bl_205 br_205 bl_out_25 br_out_25 sel_5 gnd single_level_column_mux_0
XXMUX206 bl_206 br_206 bl_out_25 br_out_25 sel_6 gnd single_level_column_mux_0
XXMUX207 bl_207 br_207 bl_out_25 br_out_25 sel_7 gnd single_level_column_mux_0
XXMUX208 bl_208 br_208 bl_out_26 br_out_26 sel_0 gnd single_level_column_mux_0
XXMUX209 bl_209 br_209 bl_out_26 br_out_26 sel_1 gnd single_level_column_mux_0
XXMUX210 bl_210 br_210 bl_out_26 br_out_26 sel_2 gnd single_level_column_mux_0
XXMUX211 bl_211 br_211 bl_out_26 br_out_26 sel_3 gnd single_level_column_mux_0
XXMUX212 bl_212 br_212 bl_out_26 br_out_26 sel_4 gnd single_level_column_mux_0
XXMUX213 bl_213 br_213 bl_out_26 br_out_26 sel_5 gnd single_level_column_mux_0
XXMUX214 bl_214 br_214 bl_out_26 br_out_26 sel_6 gnd single_level_column_mux_0
XXMUX215 bl_215 br_215 bl_out_26 br_out_26 sel_7 gnd single_level_column_mux_0
XXMUX216 bl_216 br_216 bl_out_27 br_out_27 sel_0 gnd single_level_column_mux_0
XXMUX217 bl_217 br_217 bl_out_27 br_out_27 sel_1 gnd single_level_column_mux_0
XXMUX218 bl_218 br_218 bl_out_27 br_out_27 sel_2 gnd single_level_column_mux_0
XXMUX219 bl_219 br_219 bl_out_27 br_out_27 sel_3 gnd single_level_column_mux_0
XXMUX220 bl_220 br_220 bl_out_27 br_out_27 sel_4 gnd single_level_column_mux_0
XXMUX221 bl_221 br_221 bl_out_27 br_out_27 sel_5 gnd single_level_column_mux_0
XXMUX222 bl_222 br_222 bl_out_27 br_out_27 sel_6 gnd single_level_column_mux_0
XXMUX223 bl_223 br_223 bl_out_27 br_out_27 sel_7 gnd single_level_column_mux_0
XXMUX224 bl_224 br_224 bl_out_28 br_out_28 sel_0 gnd single_level_column_mux_0
XXMUX225 bl_225 br_225 bl_out_28 br_out_28 sel_1 gnd single_level_column_mux_0
XXMUX226 bl_226 br_226 bl_out_28 br_out_28 sel_2 gnd single_level_column_mux_0
XXMUX227 bl_227 br_227 bl_out_28 br_out_28 sel_3 gnd single_level_column_mux_0
XXMUX228 bl_228 br_228 bl_out_28 br_out_28 sel_4 gnd single_level_column_mux_0
XXMUX229 bl_229 br_229 bl_out_28 br_out_28 sel_5 gnd single_level_column_mux_0
XXMUX230 bl_230 br_230 bl_out_28 br_out_28 sel_6 gnd single_level_column_mux_0
XXMUX231 bl_231 br_231 bl_out_28 br_out_28 sel_7 gnd single_level_column_mux_0
XXMUX232 bl_232 br_232 bl_out_29 br_out_29 sel_0 gnd single_level_column_mux_0
XXMUX233 bl_233 br_233 bl_out_29 br_out_29 sel_1 gnd single_level_column_mux_0
XXMUX234 bl_234 br_234 bl_out_29 br_out_29 sel_2 gnd single_level_column_mux_0
XXMUX235 bl_235 br_235 bl_out_29 br_out_29 sel_3 gnd single_level_column_mux_0
XXMUX236 bl_236 br_236 bl_out_29 br_out_29 sel_4 gnd single_level_column_mux_0
XXMUX237 bl_237 br_237 bl_out_29 br_out_29 sel_5 gnd single_level_column_mux_0
XXMUX238 bl_238 br_238 bl_out_29 br_out_29 sel_6 gnd single_level_column_mux_0
XXMUX239 bl_239 br_239 bl_out_29 br_out_29 sel_7 gnd single_level_column_mux_0
XXMUX240 bl_240 br_240 bl_out_30 br_out_30 sel_0 gnd single_level_column_mux_0
XXMUX241 bl_241 br_241 bl_out_30 br_out_30 sel_1 gnd single_level_column_mux_0
XXMUX242 bl_242 br_242 bl_out_30 br_out_30 sel_2 gnd single_level_column_mux_0
XXMUX243 bl_243 br_243 bl_out_30 br_out_30 sel_3 gnd single_level_column_mux_0
XXMUX244 bl_244 br_244 bl_out_30 br_out_30 sel_4 gnd single_level_column_mux_0
XXMUX245 bl_245 br_245 bl_out_30 br_out_30 sel_5 gnd single_level_column_mux_0
XXMUX246 bl_246 br_246 bl_out_30 br_out_30 sel_6 gnd single_level_column_mux_0
XXMUX247 bl_247 br_247 bl_out_30 br_out_30 sel_7 gnd single_level_column_mux_0
XXMUX248 bl_248 br_248 bl_out_31 br_out_31 sel_0 gnd single_level_column_mux_0
XXMUX249 bl_249 br_249 bl_out_31 br_out_31 sel_1 gnd single_level_column_mux_0
XXMUX250 bl_250 br_250 bl_out_31 br_out_31 sel_2 gnd single_level_column_mux_0
XXMUX251 bl_251 br_251 bl_out_31 br_out_31 sel_3 gnd single_level_column_mux_0
XXMUX252 bl_252 br_252 bl_out_31 br_out_31 sel_4 gnd single_level_column_mux_0
XXMUX253 bl_253 br_253 bl_out_31 br_out_31 sel_5 gnd single_level_column_mux_0
XXMUX254 bl_254 br_254 bl_out_31 br_out_31 sel_6 gnd single_level_column_mux_0
XXMUX255 bl_255 br_255 bl_out_31 br_out_31 sel_7 gnd single_level_column_mux_0
.ENDS single_level_column_mux_array_0

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT write_driver_array_0 data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 data_8 data_9 data_10 data_11 data_12 data_13 data_14 data_15 data_16 data_17 data_18 data_19 data_20 data_21 data_22 data_23 data_24 data_25 data_26 data_27 data_28 data_29 data_30 data_31 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 en vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* INPUT : data_8 
* INPUT : data_9 
* INPUT : data_10 
* INPUT : data_11 
* INPUT : data_12 
* INPUT : data_13 
* INPUT : data_14 
* INPUT : data_15 
* INPUT : data_16 
* INPUT : data_17 
* INPUT : data_18 
* INPUT : data_19 
* INPUT : data_20 
* INPUT : data_21 
* INPUT : data_22 
* INPUT : data_23 
* INPUT : data_24 
* INPUT : data_25 
* INPUT : data_26 
* INPUT : data_27 
* INPUT : data_28 
* INPUT : data_29 
* INPUT : data_30 
* INPUT : data_31 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xwrite_driver0 data_0 bl_0 br_0 en vdd gnd write_driver
Xwrite_driver8 data_1 bl_1 br_1 en vdd gnd write_driver
Xwrite_driver16 data_2 bl_2 br_2 en vdd gnd write_driver
Xwrite_driver24 data_3 bl_3 br_3 en vdd gnd write_driver
Xwrite_driver32 data_4 bl_4 br_4 en vdd gnd write_driver
Xwrite_driver40 data_5 bl_5 br_5 en vdd gnd write_driver
Xwrite_driver48 data_6 bl_6 br_6 en vdd gnd write_driver
Xwrite_driver56 data_7 bl_7 br_7 en vdd gnd write_driver
Xwrite_driver64 data_8 bl_8 br_8 en vdd gnd write_driver
Xwrite_driver72 data_9 bl_9 br_9 en vdd gnd write_driver
Xwrite_driver80 data_10 bl_10 br_10 en vdd gnd write_driver
Xwrite_driver88 data_11 bl_11 br_11 en vdd gnd write_driver
Xwrite_driver96 data_12 bl_12 br_12 en vdd gnd write_driver
Xwrite_driver104 data_13 bl_13 br_13 en vdd gnd write_driver
Xwrite_driver112 data_14 bl_14 br_14 en vdd gnd write_driver
Xwrite_driver120 data_15 bl_15 br_15 en vdd gnd write_driver
Xwrite_driver128 data_16 bl_16 br_16 en vdd gnd write_driver
Xwrite_driver136 data_17 bl_17 br_17 en vdd gnd write_driver
Xwrite_driver144 data_18 bl_18 br_18 en vdd gnd write_driver
Xwrite_driver152 data_19 bl_19 br_19 en vdd gnd write_driver
Xwrite_driver160 data_20 bl_20 br_20 en vdd gnd write_driver
Xwrite_driver168 data_21 bl_21 br_21 en vdd gnd write_driver
Xwrite_driver176 data_22 bl_22 br_22 en vdd gnd write_driver
Xwrite_driver184 data_23 bl_23 br_23 en vdd gnd write_driver
Xwrite_driver192 data_24 bl_24 br_24 en vdd gnd write_driver
Xwrite_driver200 data_25 bl_25 br_25 en vdd gnd write_driver
Xwrite_driver208 data_26 bl_26 br_26 en vdd gnd write_driver
Xwrite_driver216 data_27 bl_27 br_27 en vdd gnd write_driver
Xwrite_driver224 data_28 bl_28 br_28 en vdd gnd write_driver
Xwrite_driver232 data_29 bl_29 br_29 en vdd gnd write_driver
Xwrite_driver240 data_30 bl_30 br_30 en vdd gnd write_driver
Xwrite_driver248 data_31 bl_31 br_31 en vdd gnd write_driver
.ENDS write_driver_array_0

.SUBCKT port_data_0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout_0 dout_1 dout_2 dout_3 dout_4 dout_5 dout_6 dout_7 dout_8 dout_9 dout_10 dout_11 dout_12 dout_13 dout_14 dout_15 dout_16 dout_17 dout_18 dout_19 dout_20 dout_21 dout_22 dout_23 dout_24 dout_25 dout_26 dout_27 dout_28 dout_29 dout_30 dout_31 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 s_en p_en_bar w_en vdd gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* OUTPUT: dout_8 
* OUTPUT: dout_9 
* OUTPUT: dout_10 
* OUTPUT: dout_11 
* OUTPUT: dout_12 
* OUTPUT: dout_13 
* OUTPUT: dout_14 
* OUTPUT: dout_15 
* OUTPUT: dout_16 
* OUTPUT: dout_17 
* OUTPUT: dout_18 
* OUTPUT: dout_19 
* OUTPUT: dout_20 
* OUTPUT: dout_21 
* OUTPUT: dout_22 
* OUTPUT: dout_23 
* OUTPUT: dout_24 
* OUTPUT: dout_25 
* OUTPUT: dout_26 
* OUTPUT: dout_27 
* OUTPUT: dout_28 
* OUTPUT: dout_29 
* OUTPUT: dout_30 
* OUTPUT: dout_31 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : din_8 
* INPUT : din_9 
* INPUT : din_10 
* INPUT : din_11 
* INPUT : din_12 
* INPUT : din_13 
* INPUT : din_14 
* INPUT : din_15 
* INPUT : din_16 
* INPUT : din_17 
* INPUT : din_18 
* INPUT : din_19 
* INPUT : din_20 
* INPUT : din_21 
* INPUT : din_22 
* INPUT : din_23 
* INPUT : din_24 
* INPUT : din_25 
* INPUT : din_26 
* INPUT : din_27 
* INPUT : din_28 
* INPUT : din_29 
* INPUT : din_30 
* INPUT : din_31 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : sel_2 
* INPUT : sel_3 
* INPUT : sel_4 
* INPUT : sel_5 
* INPUT : sel_6 
* INPUT : sel_7 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0 rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 p_en_bar vdd precharge_array_0
Xsense_amp_array0 dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2 br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5 bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7 dout_8 bl_out_8 br_out_8 dout_9 bl_out_9 br_out_9 dout_10 bl_out_10 br_out_10 dout_11 bl_out_11 br_out_11 dout_12 bl_out_12 br_out_12 dout_13 bl_out_13 br_out_13 dout_14 bl_out_14 br_out_14 dout_15 bl_out_15 br_out_15 dout_16 bl_out_16 br_out_16 dout_17 bl_out_17 br_out_17 dout_18 bl_out_18 br_out_18 dout_19 bl_out_19 br_out_19 dout_20 bl_out_20 br_out_20 dout_21 bl_out_21 br_out_21 dout_22 bl_out_22 br_out_22 dout_23 bl_out_23 br_out_23 dout_24 bl_out_24 br_out_24 dout_25 bl_out_25 br_out_25 dout_26 bl_out_26 br_out_26 dout_27 bl_out_27 br_out_27 dout_28 bl_out_28 br_out_28 dout_29 bl_out_29 br_out_29 dout_30 bl_out_30 br_out_30 dout_31 bl_out_31 br_out_31 s_en vdd gnd sense_amp_array_0
Xwrite_driver_array0 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 din_8 din_9 din_10 din_11 din_12 din_13 din_14 din_15 din_16 din_17 din_18 din_19 din_20 din_21 din_22 din_23 din_24 din_25 din_26 din_27 din_28 din_29 din_30 din_31 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 w_en vdd gnd write_driver_array_0
Xcolumn_mux_array0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 bl_out_8 br_out_8 bl_out_9 br_out_9 bl_out_10 br_out_10 bl_out_11 br_out_11 bl_out_12 br_out_12 bl_out_13 br_out_13 bl_out_14 br_out_14 bl_out_15 br_out_15 bl_out_16 br_out_16 bl_out_17 br_out_17 bl_out_18 br_out_18 bl_out_19 br_out_19 bl_out_20 br_out_20 bl_out_21 br_out_21 bl_out_22 br_out_22 bl_out_23 br_out_23 bl_out_24 br_out_24 bl_out_25 br_out_25 bl_out_26 br_out_26 bl_out_27 br_out_27 bl_out_28 br_out_28 bl_out_29 br_out_29 bl_out_30 br_out_30 bl_out_31 br_out_31 gnd single_level_column_mux_array_0
.ENDS port_data_0

* ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_0

* ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

.SUBCKT pnand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_0

.SUBCKT pnand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_0

.SUBCKT hierarchical_predecode2x4_0 in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
XXpre2x4_nand_0 inbar_0 inbar_1 Z_0 vdd gnd pnand2_0
XXpre2x4_nand_1 in_0 inbar_1 Z_1 vdd gnd pnand2_0
XXpre2x4_nand_2 inbar_0 in_1 Z_2 vdd gnd pnand2_0
XXpre2x4_nand_3 in_0 in_1 Z_3 vdd gnd pnand2_0
.ENDS hierarchical_predecode2x4_0

.SUBCKT hierarchical_predecode3x8_0 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_0
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_0
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_0
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_0
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_0
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_0
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_0
Xpre_nand_inv_4 Z_4 out_4 vdd gnd pinv_0
Xpre_nand_inv_5 Z_5 out_5 vdd gnd pinv_0
Xpre_nand_inv_6 Z_6 out_6 vdd gnd pinv_0
Xpre_nand_inv_7 Z_7 out_7 vdd gnd pinv_0
XXpre3x8_nand_0 inbar_0 inbar_1 inbar_2 Z_0 vdd gnd pnand3_0
XXpre3x8_nand_1 in_0 inbar_1 inbar_2 Z_1 vdd gnd pnand3_0
XXpre3x8_nand_2 inbar_0 in_1 inbar_2 Z_2 vdd gnd pnand3_0
XXpre3x8_nand_3 in_0 in_1 inbar_2 Z_3 vdd gnd pnand3_0
XXpre3x8_nand_4 inbar_0 inbar_1 in_2 Z_4 vdd gnd pnand3_0
XXpre3x8_nand_5 in_0 inbar_1 in_2 Z_5 vdd gnd pnand3_0
XXpre3x8_nand_6 inbar_0 in_1 in_2 Z_6 vdd gnd pnand3_0
XXpre3x8_nand_7 in_0 in_1 in_2 Z_7 vdd gnd pnand3_0
.ENDS hierarchical_predecode3x8_0

.SUBCKT hierarchical_decoder_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 decode_0 decode_1 decode_2 decode_3 decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10 decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17 decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24 decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31 decode_32 decode_33 decode_34 decode_35 decode_36 decode_37 decode_38 decode_39 decode_40 decode_41 decode_42 decode_43 decode_44 decode_45 decode_46 decode_47 decode_48 decode_49 decode_50 decode_51 decode_52 decode_53 decode_54 decode_55 decode_56 decode_57 decode_58 decode_59 decode_60 decode_61 decode_62 decode_63 decode_64 decode_65 decode_66 decode_67 decode_68 decode_69 decode_70 decode_71 decode_72 decode_73 decode_74 decode_75 decode_76 decode_77 decode_78 decode_79 decode_80 decode_81 decode_82 decode_83 decode_84 decode_85 decode_86 decode_87 decode_88 decode_89 decode_90 decode_91 decode_92 decode_93 decode_94 decode_95 decode_96 decode_97 decode_98 decode_99 decode_100 decode_101 decode_102 decode_103 decode_104 decode_105 decode_106 decode_107 decode_108 decode_109 decode_110 decode_111 decode_112 decode_113 decode_114 decode_115 decode_116 decode_117 decode_118 decode_119 decode_120 decode_121 decode_122 decode_123 decode_124 decode_125 decode_126 decode_127 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* OUTPUT: decode_32 
* OUTPUT: decode_33 
* OUTPUT: decode_34 
* OUTPUT: decode_35 
* OUTPUT: decode_36 
* OUTPUT: decode_37 
* OUTPUT: decode_38 
* OUTPUT: decode_39 
* OUTPUT: decode_40 
* OUTPUT: decode_41 
* OUTPUT: decode_42 
* OUTPUT: decode_43 
* OUTPUT: decode_44 
* OUTPUT: decode_45 
* OUTPUT: decode_46 
* OUTPUT: decode_47 
* OUTPUT: decode_48 
* OUTPUT: decode_49 
* OUTPUT: decode_50 
* OUTPUT: decode_51 
* OUTPUT: decode_52 
* OUTPUT: decode_53 
* OUTPUT: decode_54 
* OUTPUT: decode_55 
* OUTPUT: decode_56 
* OUTPUT: decode_57 
* OUTPUT: decode_58 
* OUTPUT: decode_59 
* OUTPUT: decode_60 
* OUTPUT: decode_61 
* OUTPUT: decode_62 
* OUTPUT: decode_63 
* OUTPUT: decode_64 
* OUTPUT: decode_65 
* OUTPUT: decode_66 
* OUTPUT: decode_67 
* OUTPUT: decode_68 
* OUTPUT: decode_69 
* OUTPUT: decode_70 
* OUTPUT: decode_71 
* OUTPUT: decode_72 
* OUTPUT: decode_73 
* OUTPUT: decode_74 
* OUTPUT: decode_75 
* OUTPUT: decode_76 
* OUTPUT: decode_77 
* OUTPUT: decode_78 
* OUTPUT: decode_79 
* OUTPUT: decode_80 
* OUTPUT: decode_81 
* OUTPUT: decode_82 
* OUTPUT: decode_83 
* OUTPUT: decode_84 
* OUTPUT: decode_85 
* OUTPUT: decode_86 
* OUTPUT: decode_87 
* OUTPUT: decode_88 
* OUTPUT: decode_89 
* OUTPUT: decode_90 
* OUTPUT: decode_91 
* OUTPUT: decode_92 
* OUTPUT: decode_93 
* OUTPUT: decode_94 
* OUTPUT: decode_95 
* OUTPUT: decode_96 
* OUTPUT: decode_97 
* OUTPUT: decode_98 
* OUTPUT: decode_99 
* OUTPUT: decode_100 
* OUTPUT: decode_101 
* OUTPUT: decode_102 
* OUTPUT: decode_103 
* OUTPUT: decode_104 
* OUTPUT: decode_105 
* OUTPUT: decode_106 
* OUTPUT: decode_107 
* OUTPUT: decode_108 
* OUTPUT: decode_109 
* OUTPUT: decode_110 
* OUTPUT: decode_111 
* OUTPUT: decode_112 
* OUTPUT: decode_113 
* OUTPUT: decode_114 
* OUTPUT: decode_115 
* OUTPUT: decode_116 
* OUTPUT: decode_117 
* OUTPUT: decode_118 
* OUTPUT: decode_119 
* OUTPUT: decode_120 
* OUTPUT: decode_121 
* OUTPUT: decode_122 
* OUTPUT: decode_123 
* OUTPUT: decode_124 
* OUTPUT: decode_125 
* OUTPUT: decode_126 
* OUTPUT: decode_127 
* POWER : vdd 
* GROUND: gnd 
Xpre_0 addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd hierarchical_predecode2x4_0
Xpre_1 addr_2 addr_3 out_4 out_5 out_6 out_7 vdd gnd hierarchical_predecode2x4_0
Xpre3x8_0 addr_4 addr_5 addr_6 out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15 vdd gnd hierarchical_predecode3x8_0
XDEC_NAND_0 out_0 out_4 out_8 Z_0 vdd gnd pnand3_0
XDEC_NAND_16 out_0 out_4 out_9 Z_16 vdd gnd pnand3_0
XDEC_NAND_32 out_0 out_4 out_10 Z_32 vdd gnd pnand3_0
XDEC_NAND_48 out_0 out_4 out_11 Z_48 vdd gnd pnand3_0
XDEC_NAND_64 out_0 out_4 out_12 Z_64 vdd gnd pnand3_0
XDEC_NAND_80 out_0 out_4 out_13 Z_80 vdd gnd pnand3_0
XDEC_NAND_96 out_0 out_4 out_14 Z_96 vdd gnd pnand3_0
XDEC_NAND_112 out_0 out_4 out_15 Z_112 vdd gnd pnand3_0
XDEC_NAND_4 out_0 out_5 out_8 Z_4 vdd gnd pnand3_0
XDEC_NAND_20 out_0 out_5 out_9 Z_20 vdd gnd pnand3_0
XDEC_NAND_36 out_0 out_5 out_10 Z_36 vdd gnd pnand3_0
XDEC_NAND_52 out_0 out_5 out_11 Z_52 vdd gnd pnand3_0
XDEC_NAND_68 out_0 out_5 out_12 Z_68 vdd gnd pnand3_0
XDEC_NAND_84 out_0 out_5 out_13 Z_84 vdd gnd pnand3_0
XDEC_NAND_100 out_0 out_5 out_14 Z_100 vdd gnd pnand3_0
XDEC_NAND_116 out_0 out_5 out_15 Z_116 vdd gnd pnand3_0
XDEC_NAND_8 out_0 out_6 out_8 Z_8 vdd gnd pnand3_0
XDEC_NAND_24 out_0 out_6 out_9 Z_24 vdd gnd pnand3_0
XDEC_NAND_40 out_0 out_6 out_10 Z_40 vdd gnd pnand3_0
XDEC_NAND_56 out_0 out_6 out_11 Z_56 vdd gnd pnand3_0
XDEC_NAND_72 out_0 out_6 out_12 Z_72 vdd gnd pnand3_0
XDEC_NAND_88 out_0 out_6 out_13 Z_88 vdd gnd pnand3_0
XDEC_NAND_104 out_0 out_6 out_14 Z_104 vdd gnd pnand3_0
XDEC_NAND_120 out_0 out_6 out_15 Z_120 vdd gnd pnand3_0
XDEC_NAND_12 out_0 out_7 out_8 Z_12 vdd gnd pnand3_0
XDEC_NAND_28 out_0 out_7 out_9 Z_28 vdd gnd pnand3_0
XDEC_NAND_44 out_0 out_7 out_10 Z_44 vdd gnd pnand3_0
XDEC_NAND_60 out_0 out_7 out_11 Z_60 vdd gnd pnand3_0
XDEC_NAND_76 out_0 out_7 out_12 Z_76 vdd gnd pnand3_0
XDEC_NAND_92 out_0 out_7 out_13 Z_92 vdd gnd pnand3_0
XDEC_NAND_108 out_0 out_7 out_14 Z_108 vdd gnd pnand3_0
XDEC_NAND_124 out_0 out_7 out_15 Z_124 vdd gnd pnand3_0
XDEC_NAND_1 out_1 out_4 out_8 Z_1 vdd gnd pnand3_0
XDEC_NAND_17 out_1 out_4 out_9 Z_17 vdd gnd pnand3_0
XDEC_NAND_33 out_1 out_4 out_10 Z_33 vdd gnd pnand3_0
XDEC_NAND_49 out_1 out_4 out_11 Z_49 vdd gnd pnand3_0
XDEC_NAND_65 out_1 out_4 out_12 Z_65 vdd gnd pnand3_0
XDEC_NAND_81 out_1 out_4 out_13 Z_81 vdd gnd pnand3_0
XDEC_NAND_97 out_1 out_4 out_14 Z_97 vdd gnd pnand3_0
XDEC_NAND_113 out_1 out_4 out_15 Z_113 vdd gnd pnand3_0
XDEC_NAND_5 out_1 out_5 out_8 Z_5 vdd gnd pnand3_0
XDEC_NAND_21 out_1 out_5 out_9 Z_21 vdd gnd pnand3_0
XDEC_NAND_37 out_1 out_5 out_10 Z_37 vdd gnd pnand3_0
XDEC_NAND_53 out_1 out_5 out_11 Z_53 vdd gnd pnand3_0
XDEC_NAND_69 out_1 out_5 out_12 Z_69 vdd gnd pnand3_0
XDEC_NAND_85 out_1 out_5 out_13 Z_85 vdd gnd pnand3_0
XDEC_NAND_101 out_1 out_5 out_14 Z_101 vdd gnd pnand3_0
XDEC_NAND_117 out_1 out_5 out_15 Z_117 vdd gnd pnand3_0
XDEC_NAND_9 out_1 out_6 out_8 Z_9 vdd gnd pnand3_0
XDEC_NAND_25 out_1 out_6 out_9 Z_25 vdd gnd pnand3_0
XDEC_NAND_41 out_1 out_6 out_10 Z_41 vdd gnd pnand3_0
XDEC_NAND_57 out_1 out_6 out_11 Z_57 vdd gnd pnand3_0
XDEC_NAND_73 out_1 out_6 out_12 Z_73 vdd gnd pnand3_0
XDEC_NAND_89 out_1 out_6 out_13 Z_89 vdd gnd pnand3_0
XDEC_NAND_105 out_1 out_6 out_14 Z_105 vdd gnd pnand3_0
XDEC_NAND_121 out_1 out_6 out_15 Z_121 vdd gnd pnand3_0
XDEC_NAND_13 out_1 out_7 out_8 Z_13 vdd gnd pnand3_0
XDEC_NAND_29 out_1 out_7 out_9 Z_29 vdd gnd pnand3_0
XDEC_NAND_45 out_1 out_7 out_10 Z_45 vdd gnd pnand3_0
XDEC_NAND_61 out_1 out_7 out_11 Z_61 vdd gnd pnand3_0
XDEC_NAND_77 out_1 out_7 out_12 Z_77 vdd gnd pnand3_0
XDEC_NAND_93 out_1 out_7 out_13 Z_93 vdd gnd pnand3_0
XDEC_NAND_109 out_1 out_7 out_14 Z_109 vdd gnd pnand3_0
XDEC_NAND_125 out_1 out_7 out_15 Z_125 vdd gnd pnand3_0
XDEC_NAND_2 out_2 out_4 out_8 Z_2 vdd gnd pnand3_0
XDEC_NAND_18 out_2 out_4 out_9 Z_18 vdd gnd pnand3_0
XDEC_NAND_34 out_2 out_4 out_10 Z_34 vdd gnd pnand3_0
XDEC_NAND_50 out_2 out_4 out_11 Z_50 vdd gnd pnand3_0
XDEC_NAND_66 out_2 out_4 out_12 Z_66 vdd gnd pnand3_0
XDEC_NAND_82 out_2 out_4 out_13 Z_82 vdd gnd pnand3_0
XDEC_NAND_98 out_2 out_4 out_14 Z_98 vdd gnd pnand3_0
XDEC_NAND_114 out_2 out_4 out_15 Z_114 vdd gnd pnand3_0
XDEC_NAND_6 out_2 out_5 out_8 Z_6 vdd gnd pnand3_0
XDEC_NAND_22 out_2 out_5 out_9 Z_22 vdd gnd pnand3_0
XDEC_NAND_38 out_2 out_5 out_10 Z_38 vdd gnd pnand3_0
XDEC_NAND_54 out_2 out_5 out_11 Z_54 vdd gnd pnand3_0
XDEC_NAND_70 out_2 out_5 out_12 Z_70 vdd gnd pnand3_0
XDEC_NAND_86 out_2 out_5 out_13 Z_86 vdd gnd pnand3_0
XDEC_NAND_102 out_2 out_5 out_14 Z_102 vdd gnd pnand3_0
XDEC_NAND_118 out_2 out_5 out_15 Z_118 vdd gnd pnand3_0
XDEC_NAND_10 out_2 out_6 out_8 Z_10 vdd gnd pnand3_0
XDEC_NAND_26 out_2 out_6 out_9 Z_26 vdd gnd pnand3_0
XDEC_NAND_42 out_2 out_6 out_10 Z_42 vdd gnd pnand3_0
XDEC_NAND_58 out_2 out_6 out_11 Z_58 vdd gnd pnand3_0
XDEC_NAND_74 out_2 out_6 out_12 Z_74 vdd gnd pnand3_0
XDEC_NAND_90 out_2 out_6 out_13 Z_90 vdd gnd pnand3_0
XDEC_NAND_106 out_2 out_6 out_14 Z_106 vdd gnd pnand3_0
XDEC_NAND_122 out_2 out_6 out_15 Z_122 vdd gnd pnand3_0
XDEC_NAND_14 out_2 out_7 out_8 Z_14 vdd gnd pnand3_0
XDEC_NAND_30 out_2 out_7 out_9 Z_30 vdd gnd pnand3_0
XDEC_NAND_46 out_2 out_7 out_10 Z_46 vdd gnd pnand3_0
XDEC_NAND_62 out_2 out_7 out_11 Z_62 vdd gnd pnand3_0
XDEC_NAND_78 out_2 out_7 out_12 Z_78 vdd gnd pnand3_0
XDEC_NAND_94 out_2 out_7 out_13 Z_94 vdd gnd pnand3_0
XDEC_NAND_110 out_2 out_7 out_14 Z_110 vdd gnd pnand3_0
XDEC_NAND_126 out_2 out_7 out_15 Z_126 vdd gnd pnand3_0
XDEC_NAND_3 out_3 out_4 out_8 Z_3 vdd gnd pnand3_0
XDEC_NAND_19 out_3 out_4 out_9 Z_19 vdd gnd pnand3_0
XDEC_NAND_35 out_3 out_4 out_10 Z_35 vdd gnd pnand3_0
XDEC_NAND_51 out_3 out_4 out_11 Z_51 vdd gnd pnand3_0
XDEC_NAND_67 out_3 out_4 out_12 Z_67 vdd gnd pnand3_0
XDEC_NAND_83 out_3 out_4 out_13 Z_83 vdd gnd pnand3_0
XDEC_NAND_99 out_3 out_4 out_14 Z_99 vdd gnd pnand3_0
XDEC_NAND_115 out_3 out_4 out_15 Z_115 vdd gnd pnand3_0
XDEC_NAND_7 out_3 out_5 out_8 Z_7 vdd gnd pnand3_0
XDEC_NAND_23 out_3 out_5 out_9 Z_23 vdd gnd pnand3_0
XDEC_NAND_39 out_3 out_5 out_10 Z_39 vdd gnd pnand3_0
XDEC_NAND_55 out_3 out_5 out_11 Z_55 vdd gnd pnand3_0
XDEC_NAND_71 out_3 out_5 out_12 Z_71 vdd gnd pnand3_0
XDEC_NAND_87 out_3 out_5 out_13 Z_87 vdd gnd pnand3_0
XDEC_NAND_103 out_3 out_5 out_14 Z_103 vdd gnd pnand3_0
XDEC_NAND_119 out_3 out_5 out_15 Z_119 vdd gnd pnand3_0
XDEC_NAND_11 out_3 out_6 out_8 Z_11 vdd gnd pnand3_0
XDEC_NAND_27 out_3 out_6 out_9 Z_27 vdd gnd pnand3_0
XDEC_NAND_43 out_3 out_6 out_10 Z_43 vdd gnd pnand3_0
XDEC_NAND_59 out_3 out_6 out_11 Z_59 vdd gnd pnand3_0
XDEC_NAND_75 out_3 out_6 out_12 Z_75 vdd gnd pnand3_0
XDEC_NAND_91 out_3 out_6 out_13 Z_91 vdd gnd pnand3_0
XDEC_NAND_107 out_3 out_6 out_14 Z_107 vdd gnd pnand3_0
XDEC_NAND_123 out_3 out_6 out_15 Z_123 vdd gnd pnand3_0
XDEC_NAND_15 out_3 out_7 out_8 Z_15 vdd gnd pnand3_0
XDEC_NAND_31 out_3 out_7 out_9 Z_31 vdd gnd pnand3_0
XDEC_NAND_47 out_3 out_7 out_10 Z_47 vdd gnd pnand3_0
XDEC_NAND_63 out_3 out_7 out_11 Z_63 vdd gnd pnand3_0
XDEC_NAND_79 out_3 out_7 out_12 Z_79 vdd gnd pnand3_0
XDEC_NAND_95 out_3 out_7 out_13 Z_95 vdd gnd pnand3_0
XDEC_NAND_111 out_3 out_7 out_14 Z_111 vdd gnd pnand3_0
XDEC_NAND_127 out_3 out_7 out_15 Z_127 vdd gnd pnand3_0
XDEC_INV_0 Z_0 decode_0 vdd gnd pinv_0
XDEC_INV_1 Z_1 decode_1 vdd gnd pinv_0
XDEC_INV_2 Z_2 decode_2 vdd gnd pinv_0
XDEC_INV_3 Z_3 decode_3 vdd gnd pinv_0
XDEC_INV_4 Z_4 decode_4 vdd gnd pinv_0
XDEC_INV_5 Z_5 decode_5 vdd gnd pinv_0
XDEC_INV_6 Z_6 decode_6 vdd gnd pinv_0
XDEC_INV_7 Z_7 decode_7 vdd gnd pinv_0
XDEC_INV_8 Z_8 decode_8 vdd gnd pinv_0
XDEC_INV_9 Z_9 decode_9 vdd gnd pinv_0
XDEC_INV_10 Z_10 decode_10 vdd gnd pinv_0
XDEC_INV_11 Z_11 decode_11 vdd gnd pinv_0
XDEC_INV_12 Z_12 decode_12 vdd gnd pinv_0
XDEC_INV_13 Z_13 decode_13 vdd gnd pinv_0
XDEC_INV_14 Z_14 decode_14 vdd gnd pinv_0
XDEC_INV_15 Z_15 decode_15 vdd gnd pinv_0
XDEC_INV_16 Z_16 decode_16 vdd gnd pinv_0
XDEC_INV_17 Z_17 decode_17 vdd gnd pinv_0
XDEC_INV_18 Z_18 decode_18 vdd gnd pinv_0
XDEC_INV_19 Z_19 decode_19 vdd gnd pinv_0
XDEC_INV_20 Z_20 decode_20 vdd gnd pinv_0
XDEC_INV_21 Z_21 decode_21 vdd gnd pinv_0
XDEC_INV_22 Z_22 decode_22 vdd gnd pinv_0
XDEC_INV_23 Z_23 decode_23 vdd gnd pinv_0
XDEC_INV_24 Z_24 decode_24 vdd gnd pinv_0
XDEC_INV_25 Z_25 decode_25 vdd gnd pinv_0
XDEC_INV_26 Z_26 decode_26 vdd gnd pinv_0
XDEC_INV_27 Z_27 decode_27 vdd gnd pinv_0
XDEC_INV_28 Z_28 decode_28 vdd gnd pinv_0
XDEC_INV_29 Z_29 decode_29 vdd gnd pinv_0
XDEC_INV_30 Z_30 decode_30 vdd gnd pinv_0
XDEC_INV_31 Z_31 decode_31 vdd gnd pinv_0
XDEC_INV_32 Z_32 decode_32 vdd gnd pinv_0
XDEC_INV_33 Z_33 decode_33 vdd gnd pinv_0
XDEC_INV_34 Z_34 decode_34 vdd gnd pinv_0
XDEC_INV_35 Z_35 decode_35 vdd gnd pinv_0
XDEC_INV_36 Z_36 decode_36 vdd gnd pinv_0
XDEC_INV_37 Z_37 decode_37 vdd gnd pinv_0
XDEC_INV_38 Z_38 decode_38 vdd gnd pinv_0
XDEC_INV_39 Z_39 decode_39 vdd gnd pinv_0
XDEC_INV_40 Z_40 decode_40 vdd gnd pinv_0
XDEC_INV_41 Z_41 decode_41 vdd gnd pinv_0
XDEC_INV_42 Z_42 decode_42 vdd gnd pinv_0
XDEC_INV_43 Z_43 decode_43 vdd gnd pinv_0
XDEC_INV_44 Z_44 decode_44 vdd gnd pinv_0
XDEC_INV_45 Z_45 decode_45 vdd gnd pinv_0
XDEC_INV_46 Z_46 decode_46 vdd gnd pinv_0
XDEC_INV_47 Z_47 decode_47 vdd gnd pinv_0
XDEC_INV_48 Z_48 decode_48 vdd gnd pinv_0
XDEC_INV_49 Z_49 decode_49 vdd gnd pinv_0
XDEC_INV_50 Z_50 decode_50 vdd gnd pinv_0
XDEC_INV_51 Z_51 decode_51 vdd gnd pinv_0
XDEC_INV_52 Z_52 decode_52 vdd gnd pinv_0
XDEC_INV_53 Z_53 decode_53 vdd gnd pinv_0
XDEC_INV_54 Z_54 decode_54 vdd gnd pinv_0
XDEC_INV_55 Z_55 decode_55 vdd gnd pinv_0
XDEC_INV_56 Z_56 decode_56 vdd gnd pinv_0
XDEC_INV_57 Z_57 decode_57 vdd gnd pinv_0
XDEC_INV_58 Z_58 decode_58 vdd gnd pinv_0
XDEC_INV_59 Z_59 decode_59 vdd gnd pinv_0
XDEC_INV_60 Z_60 decode_60 vdd gnd pinv_0
XDEC_INV_61 Z_61 decode_61 vdd gnd pinv_0
XDEC_INV_62 Z_62 decode_62 vdd gnd pinv_0
XDEC_INV_63 Z_63 decode_63 vdd gnd pinv_0
XDEC_INV_64 Z_64 decode_64 vdd gnd pinv_0
XDEC_INV_65 Z_65 decode_65 vdd gnd pinv_0
XDEC_INV_66 Z_66 decode_66 vdd gnd pinv_0
XDEC_INV_67 Z_67 decode_67 vdd gnd pinv_0
XDEC_INV_68 Z_68 decode_68 vdd gnd pinv_0
XDEC_INV_69 Z_69 decode_69 vdd gnd pinv_0
XDEC_INV_70 Z_70 decode_70 vdd gnd pinv_0
XDEC_INV_71 Z_71 decode_71 vdd gnd pinv_0
XDEC_INV_72 Z_72 decode_72 vdd gnd pinv_0
XDEC_INV_73 Z_73 decode_73 vdd gnd pinv_0
XDEC_INV_74 Z_74 decode_74 vdd gnd pinv_0
XDEC_INV_75 Z_75 decode_75 vdd gnd pinv_0
XDEC_INV_76 Z_76 decode_76 vdd gnd pinv_0
XDEC_INV_77 Z_77 decode_77 vdd gnd pinv_0
XDEC_INV_78 Z_78 decode_78 vdd gnd pinv_0
XDEC_INV_79 Z_79 decode_79 vdd gnd pinv_0
XDEC_INV_80 Z_80 decode_80 vdd gnd pinv_0
XDEC_INV_81 Z_81 decode_81 vdd gnd pinv_0
XDEC_INV_82 Z_82 decode_82 vdd gnd pinv_0
XDEC_INV_83 Z_83 decode_83 vdd gnd pinv_0
XDEC_INV_84 Z_84 decode_84 vdd gnd pinv_0
XDEC_INV_85 Z_85 decode_85 vdd gnd pinv_0
XDEC_INV_86 Z_86 decode_86 vdd gnd pinv_0
XDEC_INV_87 Z_87 decode_87 vdd gnd pinv_0
XDEC_INV_88 Z_88 decode_88 vdd gnd pinv_0
XDEC_INV_89 Z_89 decode_89 vdd gnd pinv_0
XDEC_INV_90 Z_90 decode_90 vdd gnd pinv_0
XDEC_INV_91 Z_91 decode_91 vdd gnd pinv_0
XDEC_INV_92 Z_92 decode_92 vdd gnd pinv_0
XDEC_INV_93 Z_93 decode_93 vdd gnd pinv_0
XDEC_INV_94 Z_94 decode_94 vdd gnd pinv_0
XDEC_INV_95 Z_95 decode_95 vdd gnd pinv_0
XDEC_INV_96 Z_96 decode_96 vdd gnd pinv_0
XDEC_INV_97 Z_97 decode_97 vdd gnd pinv_0
XDEC_INV_98 Z_98 decode_98 vdd gnd pinv_0
XDEC_INV_99 Z_99 decode_99 vdd gnd pinv_0
XDEC_INV_100 Z_100 decode_100 vdd gnd pinv_0
XDEC_INV_101 Z_101 decode_101 vdd gnd pinv_0
XDEC_INV_102 Z_102 decode_102 vdd gnd pinv_0
XDEC_INV_103 Z_103 decode_103 vdd gnd pinv_0
XDEC_INV_104 Z_104 decode_104 vdd gnd pinv_0
XDEC_INV_105 Z_105 decode_105 vdd gnd pinv_0
XDEC_INV_106 Z_106 decode_106 vdd gnd pinv_0
XDEC_INV_107 Z_107 decode_107 vdd gnd pinv_0
XDEC_INV_108 Z_108 decode_108 vdd gnd pinv_0
XDEC_INV_109 Z_109 decode_109 vdd gnd pinv_0
XDEC_INV_110 Z_110 decode_110 vdd gnd pinv_0
XDEC_INV_111 Z_111 decode_111 vdd gnd pinv_0
XDEC_INV_112 Z_112 decode_112 vdd gnd pinv_0
XDEC_INV_113 Z_113 decode_113 vdd gnd pinv_0
XDEC_INV_114 Z_114 decode_114 vdd gnd pinv_0
XDEC_INV_115 Z_115 decode_115 vdd gnd pinv_0
XDEC_INV_116 Z_116 decode_116 vdd gnd pinv_0
XDEC_INV_117 Z_117 decode_117 vdd gnd pinv_0
XDEC_INV_118 Z_118 decode_118 vdd gnd pinv_0
XDEC_INV_119 Z_119 decode_119 vdd gnd pinv_0
XDEC_INV_120 Z_120 decode_120 vdd gnd pinv_0
XDEC_INV_121 Z_121 decode_121 vdd gnd pinv_0
XDEC_INV_122 Z_122 decode_122 vdd gnd pinv_0
XDEC_INV_123 Z_123 decode_123 vdd gnd pinv_0
XDEC_INV_124 Z_124 decode_124 vdd gnd pinv_0
XDEC_INV_125 Z_125 decode_125 vdd gnd pinv_0
XDEC_INV_126 Z_126 decode_126 vdd gnd pinv_0
XDEC_INV_127 Z_127 decode_127 vdd gnd pinv_0
.ENDS hierarchical_decoder_0

.SUBCKT pinv_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_1

* ptx M{0} {1} nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_2

* ptx M{0} {1} nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

.SUBCKT pinv_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_3

* ptx M{0} {1} nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

.SUBCKT pinv_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.0925u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_4

* ptx M{0} {1} nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p

* ptx M{0} {1} pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p

.SUBCKT pinv_5 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=80 w=0.28750000000000003u l=0.05u pd=0.68u ps=0.68u as=0.04p ad=0.04p
Mpinv_nmos Z A gnd gnd nmos_vtg m=80 w=0.095u l=0.05u pd=0.29u ps=0.29u as=0.01p ad=0.01p
.ENDS pinv_5

.SUBCKT pdriver_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_1
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_1
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_1
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_2
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_3
Xbuf_inv6 Zb5_int Zb6_int vdd gnd pinv_4
Xbuf_inv7 Zb6_int Z vdd gnd pinv_5
.ENDS pdriver_0

.SUBCKT wordline_driver_0 in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12 in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23 in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34 in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45 in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56 in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67 in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78 in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89 in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100 in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110 in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120 in_121 in_122 in_123 in_124 in_125 in_126 in_127 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
Xwl_driver_nand0 en in_0 wl_bar_0 vdd gnd pnand2_0
Xwl_driver_inv0 wl_bar_0 wl_0 vdd gnd pdriver_0
Xwl_driver_nand1 en in_1 wl_bar_1 vdd gnd pnand2_0
Xwl_driver_inv1 wl_bar_1 wl_1 vdd gnd pdriver_0
Xwl_driver_nand2 en in_2 wl_bar_2 vdd gnd pnand2_0
Xwl_driver_inv2 wl_bar_2 wl_2 vdd gnd pdriver_0
Xwl_driver_nand3 en in_3 wl_bar_3 vdd gnd pnand2_0
Xwl_driver_inv3 wl_bar_3 wl_3 vdd gnd pdriver_0
Xwl_driver_nand4 en in_4 wl_bar_4 vdd gnd pnand2_0
Xwl_driver_inv4 wl_bar_4 wl_4 vdd gnd pdriver_0
Xwl_driver_nand5 en in_5 wl_bar_5 vdd gnd pnand2_0
Xwl_driver_inv5 wl_bar_5 wl_5 vdd gnd pdriver_0
Xwl_driver_nand6 en in_6 wl_bar_6 vdd gnd pnand2_0
Xwl_driver_inv6 wl_bar_6 wl_6 vdd gnd pdriver_0
Xwl_driver_nand7 en in_7 wl_bar_7 vdd gnd pnand2_0
Xwl_driver_inv7 wl_bar_7 wl_7 vdd gnd pdriver_0
Xwl_driver_nand8 en in_8 wl_bar_8 vdd gnd pnand2_0
Xwl_driver_inv8 wl_bar_8 wl_8 vdd gnd pdriver_0
Xwl_driver_nand9 en in_9 wl_bar_9 vdd gnd pnand2_0
Xwl_driver_inv9 wl_bar_9 wl_9 vdd gnd pdriver_0
Xwl_driver_nand10 en in_10 wl_bar_10 vdd gnd pnand2_0
Xwl_driver_inv10 wl_bar_10 wl_10 vdd gnd pdriver_0
Xwl_driver_nand11 en in_11 wl_bar_11 vdd gnd pnand2_0
Xwl_driver_inv11 wl_bar_11 wl_11 vdd gnd pdriver_0
Xwl_driver_nand12 en in_12 wl_bar_12 vdd gnd pnand2_0
Xwl_driver_inv12 wl_bar_12 wl_12 vdd gnd pdriver_0
Xwl_driver_nand13 en in_13 wl_bar_13 vdd gnd pnand2_0
Xwl_driver_inv13 wl_bar_13 wl_13 vdd gnd pdriver_0
Xwl_driver_nand14 en in_14 wl_bar_14 vdd gnd pnand2_0
Xwl_driver_inv14 wl_bar_14 wl_14 vdd gnd pdriver_0
Xwl_driver_nand15 en in_15 wl_bar_15 vdd gnd pnand2_0
Xwl_driver_inv15 wl_bar_15 wl_15 vdd gnd pdriver_0
Xwl_driver_nand16 en in_16 wl_bar_16 vdd gnd pnand2_0
Xwl_driver_inv16 wl_bar_16 wl_16 vdd gnd pdriver_0
Xwl_driver_nand17 en in_17 wl_bar_17 vdd gnd pnand2_0
Xwl_driver_inv17 wl_bar_17 wl_17 vdd gnd pdriver_0
Xwl_driver_nand18 en in_18 wl_bar_18 vdd gnd pnand2_0
Xwl_driver_inv18 wl_bar_18 wl_18 vdd gnd pdriver_0
Xwl_driver_nand19 en in_19 wl_bar_19 vdd gnd pnand2_0
Xwl_driver_inv19 wl_bar_19 wl_19 vdd gnd pdriver_0
Xwl_driver_nand20 en in_20 wl_bar_20 vdd gnd pnand2_0
Xwl_driver_inv20 wl_bar_20 wl_20 vdd gnd pdriver_0
Xwl_driver_nand21 en in_21 wl_bar_21 vdd gnd pnand2_0
Xwl_driver_inv21 wl_bar_21 wl_21 vdd gnd pdriver_0
Xwl_driver_nand22 en in_22 wl_bar_22 vdd gnd pnand2_0
Xwl_driver_inv22 wl_bar_22 wl_22 vdd gnd pdriver_0
Xwl_driver_nand23 en in_23 wl_bar_23 vdd gnd pnand2_0
Xwl_driver_inv23 wl_bar_23 wl_23 vdd gnd pdriver_0
Xwl_driver_nand24 en in_24 wl_bar_24 vdd gnd pnand2_0
Xwl_driver_inv24 wl_bar_24 wl_24 vdd gnd pdriver_0
Xwl_driver_nand25 en in_25 wl_bar_25 vdd gnd pnand2_0
Xwl_driver_inv25 wl_bar_25 wl_25 vdd gnd pdriver_0
Xwl_driver_nand26 en in_26 wl_bar_26 vdd gnd pnand2_0
Xwl_driver_inv26 wl_bar_26 wl_26 vdd gnd pdriver_0
Xwl_driver_nand27 en in_27 wl_bar_27 vdd gnd pnand2_0
Xwl_driver_inv27 wl_bar_27 wl_27 vdd gnd pdriver_0
Xwl_driver_nand28 en in_28 wl_bar_28 vdd gnd pnand2_0
Xwl_driver_inv28 wl_bar_28 wl_28 vdd gnd pdriver_0
Xwl_driver_nand29 en in_29 wl_bar_29 vdd gnd pnand2_0
Xwl_driver_inv29 wl_bar_29 wl_29 vdd gnd pdriver_0
Xwl_driver_nand30 en in_30 wl_bar_30 vdd gnd pnand2_0
Xwl_driver_inv30 wl_bar_30 wl_30 vdd gnd pdriver_0
Xwl_driver_nand31 en in_31 wl_bar_31 vdd gnd pnand2_0
Xwl_driver_inv31 wl_bar_31 wl_31 vdd gnd pdriver_0
Xwl_driver_nand32 en in_32 wl_bar_32 vdd gnd pnand2_0
Xwl_driver_inv32 wl_bar_32 wl_32 vdd gnd pdriver_0
Xwl_driver_nand33 en in_33 wl_bar_33 vdd gnd pnand2_0
Xwl_driver_inv33 wl_bar_33 wl_33 vdd gnd pdriver_0
Xwl_driver_nand34 en in_34 wl_bar_34 vdd gnd pnand2_0
Xwl_driver_inv34 wl_bar_34 wl_34 vdd gnd pdriver_0
Xwl_driver_nand35 en in_35 wl_bar_35 vdd gnd pnand2_0
Xwl_driver_inv35 wl_bar_35 wl_35 vdd gnd pdriver_0
Xwl_driver_nand36 en in_36 wl_bar_36 vdd gnd pnand2_0
Xwl_driver_inv36 wl_bar_36 wl_36 vdd gnd pdriver_0
Xwl_driver_nand37 en in_37 wl_bar_37 vdd gnd pnand2_0
Xwl_driver_inv37 wl_bar_37 wl_37 vdd gnd pdriver_0
Xwl_driver_nand38 en in_38 wl_bar_38 vdd gnd pnand2_0
Xwl_driver_inv38 wl_bar_38 wl_38 vdd gnd pdriver_0
Xwl_driver_nand39 en in_39 wl_bar_39 vdd gnd pnand2_0
Xwl_driver_inv39 wl_bar_39 wl_39 vdd gnd pdriver_0
Xwl_driver_nand40 en in_40 wl_bar_40 vdd gnd pnand2_0
Xwl_driver_inv40 wl_bar_40 wl_40 vdd gnd pdriver_0
Xwl_driver_nand41 en in_41 wl_bar_41 vdd gnd pnand2_0
Xwl_driver_inv41 wl_bar_41 wl_41 vdd gnd pdriver_0
Xwl_driver_nand42 en in_42 wl_bar_42 vdd gnd pnand2_0
Xwl_driver_inv42 wl_bar_42 wl_42 vdd gnd pdriver_0
Xwl_driver_nand43 en in_43 wl_bar_43 vdd gnd pnand2_0
Xwl_driver_inv43 wl_bar_43 wl_43 vdd gnd pdriver_0
Xwl_driver_nand44 en in_44 wl_bar_44 vdd gnd pnand2_0
Xwl_driver_inv44 wl_bar_44 wl_44 vdd gnd pdriver_0
Xwl_driver_nand45 en in_45 wl_bar_45 vdd gnd pnand2_0
Xwl_driver_inv45 wl_bar_45 wl_45 vdd gnd pdriver_0
Xwl_driver_nand46 en in_46 wl_bar_46 vdd gnd pnand2_0
Xwl_driver_inv46 wl_bar_46 wl_46 vdd gnd pdriver_0
Xwl_driver_nand47 en in_47 wl_bar_47 vdd gnd pnand2_0
Xwl_driver_inv47 wl_bar_47 wl_47 vdd gnd pdriver_0
Xwl_driver_nand48 en in_48 wl_bar_48 vdd gnd pnand2_0
Xwl_driver_inv48 wl_bar_48 wl_48 vdd gnd pdriver_0
Xwl_driver_nand49 en in_49 wl_bar_49 vdd gnd pnand2_0
Xwl_driver_inv49 wl_bar_49 wl_49 vdd gnd pdriver_0
Xwl_driver_nand50 en in_50 wl_bar_50 vdd gnd pnand2_0
Xwl_driver_inv50 wl_bar_50 wl_50 vdd gnd pdriver_0
Xwl_driver_nand51 en in_51 wl_bar_51 vdd gnd pnand2_0
Xwl_driver_inv51 wl_bar_51 wl_51 vdd gnd pdriver_0
Xwl_driver_nand52 en in_52 wl_bar_52 vdd gnd pnand2_0
Xwl_driver_inv52 wl_bar_52 wl_52 vdd gnd pdriver_0
Xwl_driver_nand53 en in_53 wl_bar_53 vdd gnd pnand2_0
Xwl_driver_inv53 wl_bar_53 wl_53 vdd gnd pdriver_0
Xwl_driver_nand54 en in_54 wl_bar_54 vdd gnd pnand2_0
Xwl_driver_inv54 wl_bar_54 wl_54 vdd gnd pdriver_0
Xwl_driver_nand55 en in_55 wl_bar_55 vdd gnd pnand2_0
Xwl_driver_inv55 wl_bar_55 wl_55 vdd gnd pdriver_0
Xwl_driver_nand56 en in_56 wl_bar_56 vdd gnd pnand2_0
Xwl_driver_inv56 wl_bar_56 wl_56 vdd gnd pdriver_0
Xwl_driver_nand57 en in_57 wl_bar_57 vdd gnd pnand2_0
Xwl_driver_inv57 wl_bar_57 wl_57 vdd gnd pdriver_0
Xwl_driver_nand58 en in_58 wl_bar_58 vdd gnd pnand2_0
Xwl_driver_inv58 wl_bar_58 wl_58 vdd gnd pdriver_0
Xwl_driver_nand59 en in_59 wl_bar_59 vdd gnd pnand2_0
Xwl_driver_inv59 wl_bar_59 wl_59 vdd gnd pdriver_0
Xwl_driver_nand60 en in_60 wl_bar_60 vdd gnd pnand2_0
Xwl_driver_inv60 wl_bar_60 wl_60 vdd gnd pdriver_0
Xwl_driver_nand61 en in_61 wl_bar_61 vdd gnd pnand2_0
Xwl_driver_inv61 wl_bar_61 wl_61 vdd gnd pdriver_0
Xwl_driver_nand62 en in_62 wl_bar_62 vdd gnd pnand2_0
Xwl_driver_inv62 wl_bar_62 wl_62 vdd gnd pdriver_0
Xwl_driver_nand63 en in_63 wl_bar_63 vdd gnd pnand2_0
Xwl_driver_inv63 wl_bar_63 wl_63 vdd gnd pdriver_0
Xwl_driver_nand64 en in_64 wl_bar_64 vdd gnd pnand2_0
Xwl_driver_inv64 wl_bar_64 wl_64 vdd gnd pdriver_0
Xwl_driver_nand65 en in_65 wl_bar_65 vdd gnd pnand2_0
Xwl_driver_inv65 wl_bar_65 wl_65 vdd gnd pdriver_0
Xwl_driver_nand66 en in_66 wl_bar_66 vdd gnd pnand2_0
Xwl_driver_inv66 wl_bar_66 wl_66 vdd gnd pdriver_0
Xwl_driver_nand67 en in_67 wl_bar_67 vdd gnd pnand2_0
Xwl_driver_inv67 wl_bar_67 wl_67 vdd gnd pdriver_0
Xwl_driver_nand68 en in_68 wl_bar_68 vdd gnd pnand2_0
Xwl_driver_inv68 wl_bar_68 wl_68 vdd gnd pdriver_0
Xwl_driver_nand69 en in_69 wl_bar_69 vdd gnd pnand2_0
Xwl_driver_inv69 wl_bar_69 wl_69 vdd gnd pdriver_0
Xwl_driver_nand70 en in_70 wl_bar_70 vdd gnd pnand2_0
Xwl_driver_inv70 wl_bar_70 wl_70 vdd gnd pdriver_0
Xwl_driver_nand71 en in_71 wl_bar_71 vdd gnd pnand2_0
Xwl_driver_inv71 wl_bar_71 wl_71 vdd gnd pdriver_0
Xwl_driver_nand72 en in_72 wl_bar_72 vdd gnd pnand2_0
Xwl_driver_inv72 wl_bar_72 wl_72 vdd gnd pdriver_0
Xwl_driver_nand73 en in_73 wl_bar_73 vdd gnd pnand2_0
Xwl_driver_inv73 wl_bar_73 wl_73 vdd gnd pdriver_0
Xwl_driver_nand74 en in_74 wl_bar_74 vdd gnd pnand2_0
Xwl_driver_inv74 wl_bar_74 wl_74 vdd gnd pdriver_0
Xwl_driver_nand75 en in_75 wl_bar_75 vdd gnd pnand2_0
Xwl_driver_inv75 wl_bar_75 wl_75 vdd gnd pdriver_0
Xwl_driver_nand76 en in_76 wl_bar_76 vdd gnd pnand2_0
Xwl_driver_inv76 wl_bar_76 wl_76 vdd gnd pdriver_0
Xwl_driver_nand77 en in_77 wl_bar_77 vdd gnd pnand2_0
Xwl_driver_inv77 wl_bar_77 wl_77 vdd gnd pdriver_0
Xwl_driver_nand78 en in_78 wl_bar_78 vdd gnd pnand2_0
Xwl_driver_inv78 wl_bar_78 wl_78 vdd gnd pdriver_0
Xwl_driver_nand79 en in_79 wl_bar_79 vdd gnd pnand2_0
Xwl_driver_inv79 wl_bar_79 wl_79 vdd gnd pdriver_0
Xwl_driver_nand80 en in_80 wl_bar_80 vdd gnd pnand2_0
Xwl_driver_inv80 wl_bar_80 wl_80 vdd gnd pdriver_0
Xwl_driver_nand81 en in_81 wl_bar_81 vdd gnd pnand2_0
Xwl_driver_inv81 wl_bar_81 wl_81 vdd gnd pdriver_0
Xwl_driver_nand82 en in_82 wl_bar_82 vdd gnd pnand2_0
Xwl_driver_inv82 wl_bar_82 wl_82 vdd gnd pdriver_0
Xwl_driver_nand83 en in_83 wl_bar_83 vdd gnd pnand2_0
Xwl_driver_inv83 wl_bar_83 wl_83 vdd gnd pdriver_0
Xwl_driver_nand84 en in_84 wl_bar_84 vdd gnd pnand2_0
Xwl_driver_inv84 wl_bar_84 wl_84 vdd gnd pdriver_0
Xwl_driver_nand85 en in_85 wl_bar_85 vdd gnd pnand2_0
Xwl_driver_inv85 wl_bar_85 wl_85 vdd gnd pdriver_0
Xwl_driver_nand86 en in_86 wl_bar_86 vdd gnd pnand2_0
Xwl_driver_inv86 wl_bar_86 wl_86 vdd gnd pdriver_0
Xwl_driver_nand87 en in_87 wl_bar_87 vdd gnd pnand2_0
Xwl_driver_inv87 wl_bar_87 wl_87 vdd gnd pdriver_0
Xwl_driver_nand88 en in_88 wl_bar_88 vdd gnd pnand2_0
Xwl_driver_inv88 wl_bar_88 wl_88 vdd gnd pdriver_0
Xwl_driver_nand89 en in_89 wl_bar_89 vdd gnd pnand2_0
Xwl_driver_inv89 wl_bar_89 wl_89 vdd gnd pdriver_0
Xwl_driver_nand90 en in_90 wl_bar_90 vdd gnd pnand2_0
Xwl_driver_inv90 wl_bar_90 wl_90 vdd gnd pdriver_0
Xwl_driver_nand91 en in_91 wl_bar_91 vdd gnd pnand2_0
Xwl_driver_inv91 wl_bar_91 wl_91 vdd gnd pdriver_0
Xwl_driver_nand92 en in_92 wl_bar_92 vdd gnd pnand2_0
Xwl_driver_inv92 wl_bar_92 wl_92 vdd gnd pdriver_0
Xwl_driver_nand93 en in_93 wl_bar_93 vdd gnd pnand2_0
Xwl_driver_inv93 wl_bar_93 wl_93 vdd gnd pdriver_0
Xwl_driver_nand94 en in_94 wl_bar_94 vdd gnd pnand2_0
Xwl_driver_inv94 wl_bar_94 wl_94 vdd gnd pdriver_0
Xwl_driver_nand95 en in_95 wl_bar_95 vdd gnd pnand2_0
Xwl_driver_inv95 wl_bar_95 wl_95 vdd gnd pdriver_0
Xwl_driver_nand96 en in_96 wl_bar_96 vdd gnd pnand2_0
Xwl_driver_inv96 wl_bar_96 wl_96 vdd gnd pdriver_0
Xwl_driver_nand97 en in_97 wl_bar_97 vdd gnd pnand2_0
Xwl_driver_inv97 wl_bar_97 wl_97 vdd gnd pdriver_0
Xwl_driver_nand98 en in_98 wl_bar_98 vdd gnd pnand2_0
Xwl_driver_inv98 wl_bar_98 wl_98 vdd gnd pdriver_0
Xwl_driver_nand99 en in_99 wl_bar_99 vdd gnd pnand2_0
Xwl_driver_inv99 wl_bar_99 wl_99 vdd gnd pdriver_0
Xwl_driver_nand100 en in_100 wl_bar_100 vdd gnd pnand2_0
Xwl_driver_inv100 wl_bar_100 wl_100 vdd gnd pdriver_0
Xwl_driver_nand101 en in_101 wl_bar_101 vdd gnd pnand2_0
Xwl_driver_inv101 wl_bar_101 wl_101 vdd gnd pdriver_0
Xwl_driver_nand102 en in_102 wl_bar_102 vdd gnd pnand2_0
Xwl_driver_inv102 wl_bar_102 wl_102 vdd gnd pdriver_0
Xwl_driver_nand103 en in_103 wl_bar_103 vdd gnd pnand2_0
Xwl_driver_inv103 wl_bar_103 wl_103 vdd gnd pdriver_0
Xwl_driver_nand104 en in_104 wl_bar_104 vdd gnd pnand2_0
Xwl_driver_inv104 wl_bar_104 wl_104 vdd gnd pdriver_0
Xwl_driver_nand105 en in_105 wl_bar_105 vdd gnd pnand2_0
Xwl_driver_inv105 wl_bar_105 wl_105 vdd gnd pdriver_0
Xwl_driver_nand106 en in_106 wl_bar_106 vdd gnd pnand2_0
Xwl_driver_inv106 wl_bar_106 wl_106 vdd gnd pdriver_0
Xwl_driver_nand107 en in_107 wl_bar_107 vdd gnd pnand2_0
Xwl_driver_inv107 wl_bar_107 wl_107 vdd gnd pdriver_0
Xwl_driver_nand108 en in_108 wl_bar_108 vdd gnd pnand2_0
Xwl_driver_inv108 wl_bar_108 wl_108 vdd gnd pdriver_0
Xwl_driver_nand109 en in_109 wl_bar_109 vdd gnd pnand2_0
Xwl_driver_inv109 wl_bar_109 wl_109 vdd gnd pdriver_0
Xwl_driver_nand110 en in_110 wl_bar_110 vdd gnd pnand2_0
Xwl_driver_inv110 wl_bar_110 wl_110 vdd gnd pdriver_0
Xwl_driver_nand111 en in_111 wl_bar_111 vdd gnd pnand2_0
Xwl_driver_inv111 wl_bar_111 wl_111 vdd gnd pdriver_0
Xwl_driver_nand112 en in_112 wl_bar_112 vdd gnd pnand2_0
Xwl_driver_inv112 wl_bar_112 wl_112 vdd gnd pdriver_0
Xwl_driver_nand113 en in_113 wl_bar_113 vdd gnd pnand2_0
Xwl_driver_inv113 wl_bar_113 wl_113 vdd gnd pdriver_0
Xwl_driver_nand114 en in_114 wl_bar_114 vdd gnd pnand2_0
Xwl_driver_inv114 wl_bar_114 wl_114 vdd gnd pdriver_0
Xwl_driver_nand115 en in_115 wl_bar_115 vdd gnd pnand2_0
Xwl_driver_inv115 wl_bar_115 wl_115 vdd gnd pdriver_0
Xwl_driver_nand116 en in_116 wl_bar_116 vdd gnd pnand2_0
Xwl_driver_inv116 wl_bar_116 wl_116 vdd gnd pdriver_0
Xwl_driver_nand117 en in_117 wl_bar_117 vdd gnd pnand2_0
Xwl_driver_inv117 wl_bar_117 wl_117 vdd gnd pdriver_0
Xwl_driver_nand118 en in_118 wl_bar_118 vdd gnd pnand2_0
Xwl_driver_inv118 wl_bar_118 wl_118 vdd gnd pdriver_0
Xwl_driver_nand119 en in_119 wl_bar_119 vdd gnd pnand2_0
Xwl_driver_inv119 wl_bar_119 wl_119 vdd gnd pdriver_0
Xwl_driver_nand120 en in_120 wl_bar_120 vdd gnd pnand2_0
Xwl_driver_inv120 wl_bar_120 wl_120 vdd gnd pdriver_0
Xwl_driver_nand121 en in_121 wl_bar_121 vdd gnd pnand2_0
Xwl_driver_inv121 wl_bar_121 wl_121 vdd gnd pdriver_0
Xwl_driver_nand122 en in_122 wl_bar_122 vdd gnd pnand2_0
Xwl_driver_inv122 wl_bar_122 wl_122 vdd gnd pdriver_0
Xwl_driver_nand123 en in_123 wl_bar_123 vdd gnd pnand2_0
Xwl_driver_inv123 wl_bar_123 wl_123 vdd gnd pdriver_0
Xwl_driver_nand124 en in_124 wl_bar_124 vdd gnd pnand2_0
Xwl_driver_inv124 wl_bar_124 wl_124 vdd gnd pdriver_0
Xwl_driver_nand125 en in_125 wl_bar_125 vdd gnd pnand2_0
Xwl_driver_inv125 wl_bar_125 wl_125 vdd gnd pdriver_0
Xwl_driver_nand126 en in_126 wl_bar_126 vdd gnd pnand2_0
Xwl_driver_inv126 wl_bar_126 wl_126 vdd gnd pdriver_0
Xwl_driver_nand127 en in_127 wl_bar_127 vdd gnd pnand2_0
Xwl_driver_inv127 wl_bar_127 wl_127 vdd gnd pdriver_0
.ENDS wordline_driver_0

.SUBCKT port_address_0 addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* OUTPUT: wl_89 
* OUTPUT: wl_90 
* OUTPUT: wl_91 
* OUTPUT: wl_92 
* OUTPUT: wl_93 
* OUTPUT: wl_94 
* OUTPUT: wl_95 
* OUTPUT: wl_96 
* OUTPUT: wl_97 
* OUTPUT: wl_98 
* OUTPUT: wl_99 
* OUTPUT: wl_100 
* OUTPUT: wl_101 
* OUTPUT: wl_102 
* OUTPUT: wl_103 
* OUTPUT: wl_104 
* OUTPUT: wl_105 
* OUTPUT: wl_106 
* OUTPUT: wl_107 
* OUTPUT: wl_108 
* OUTPUT: wl_109 
* OUTPUT: wl_110 
* OUTPUT: wl_111 
* OUTPUT: wl_112 
* OUTPUT: wl_113 
* OUTPUT: wl_114 
* OUTPUT: wl_115 
* OUTPUT: wl_116 
* OUTPUT: wl_117 
* OUTPUT: wl_118 
* OUTPUT: wl_119 
* OUTPUT: wl_120 
* OUTPUT: wl_121 
* OUTPUT: wl_122 
* OUTPUT: wl_123 
* OUTPUT: wl_124 
* OUTPUT: wl_125 
* OUTPUT: wl_126 
* OUTPUT: wl_127 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 vdd gnd hierarchical_decoder_0
Xwordline_driver dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30 dec_out_31 dec_out_32 dec_out_33 dec_out_34 dec_out_35 dec_out_36 dec_out_37 dec_out_38 dec_out_39 dec_out_40 dec_out_41 dec_out_42 dec_out_43 dec_out_44 dec_out_45 dec_out_46 dec_out_47 dec_out_48 dec_out_49 dec_out_50 dec_out_51 dec_out_52 dec_out_53 dec_out_54 dec_out_55 dec_out_56 dec_out_57 dec_out_58 dec_out_59 dec_out_60 dec_out_61 dec_out_62 dec_out_63 dec_out_64 dec_out_65 dec_out_66 dec_out_67 dec_out_68 dec_out_69 dec_out_70 dec_out_71 dec_out_72 dec_out_73 dec_out_74 dec_out_75 dec_out_76 dec_out_77 dec_out_78 dec_out_79 dec_out_80 dec_out_81 dec_out_82 dec_out_83 dec_out_84 dec_out_85 dec_out_86 dec_out_87 dec_out_88 dec_out_89 dec_out_90 dec_out_91 dec_out_92 dec_out_93 dec_out_94 dec_out_95 dec_out_96 dec_out_97 dec_out_98 dec_out_99 dec_out_100 dec_out_101 dec_out_102 dec_out_103 dec_out_104 dec_out_105 dec_out_106 dec_out_107 dec_out_108 dec_out_109 dec_out_110 dec_out_111 dec_out_112 dec_out_113 dec_out_114 dec_out_115 dec_out_116 dec_out_117 dec_out_118 dec_out_119 dec_out_120 dec_out_121 dec_out_122 dec_out_123 dec_out_124 dec_out_125 dec_out_126 dec_out_127 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_en vdd gnd wordline_driver_0
.ENDS port_address_0

.SUBCKT cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd cell_6t
Xbit_r1_c1 bl_1 br_1 wl_1 vdd gnd cell_6t
Xbit_r2_c1 bl_1 br_1 wl_2 vdd gnd cell_6t
Xbit_r3_c1 bl_1 br_1 wl_3 vdd gnd cell_6t
Xbit_r4_c1 bl_1 br_1 wl_4 vdd gnd cell_6t
Xbit_r5_c1 bl_1 br_1 wl_5 vdd gnd cell_6t
Xbit_r6_c1 bl_1 br_1 wl_6 vdd gnd cell_6t
Xbit_r7_c1 bl_1 br_1 wl_7 vdd gnd cell_6t
Xbit_r8_c1 bl_1 br_1 wl_8 vdd gnd cell_6t
Xbit_r9_c1 bl_1 br_1 wl_9 vdd gnd cell_6t
Xbit_r10_c1 bl_1 br_1 wl_10 vdd gnd cell_6t
Xbit_r11_c1 bl_1 br_1 wl_11 vdd gnd cell_6t
Xbit_r12_c1 bl_1 br_1 wl_12 vdd gnd cell_6t
Xbit_r13_c1 bl_1 br_1 wl_13 vdd gnd cell_6t
Xbit_r14_c1 bl_1 br_1 wl_14 vdd gnd cell_6t
Xbit_r15_c1 bl_1 br_1 wl_15 vdd gnd cell_6t
Xbit_r16_c1 bl_1 br_1 wl_16 vdd gnd cell_6t
Xbit_r17_c1 bl_1 br_1 wl_17 vdd gnd cell_6t
Xbit_r18_c1 bl_1 br_1 wl_18 vdd gnd cell_6t
Xbit_r19_c1 bl_1 br_1 wl_19 vdd gnd cell_6t
Xbit_r20_c1 bl_1 br_1 wl_20 vdd gnd cell_6t
Xbit_r21_c1 bl_1 br_1 wl_21 vdd gnd cell_6t
Xbit_r22_c1 bl_1 br_1 wl_22 vdd gnd cell_6t
Xbit_r23_c1 bl_1 br_1 wl_23 vdd gnd cell_6t
Xbit_r24_c1 bl_1 br_1 wl_24 vdd gnd cell_6t
Xbit_r25_c1 bl_1 br_1 wl_25 vdd gnd cell_6t
Xbit_r26_c1 bl_1 br_1 wl_26 vdd gnd cell_6t
Xbit_r27_c1 bl_1 br_1 wl_27 vdd gnd cell_6t
Xbit_r28_c1 bl_1 br_1 wl_28 vdd gnd cell_6t
Xbit_r29_c1 bl_1 br_1 wl_29 vdd gnd cell_6t
Xbit_r30_c1 bl_1 br_1 wl_30 vdd gnd cell_6t
Xbit_r31_c1 bl_1 br_1 wl_31 vdd gnd cell_6t
Xbit_r32_c1 bl_1 br_1 wl_32 vdd gnd cell_6t
Xbit_r33_c1 bl_1 br_1 wl_33 vdd gnd cell_6t
Xbit_r34_c1 bl_1 br_1 wl_34 vdd gnd cell_6t
Xbit_r35_c1 bl_1 br_1 wl_35 vdd gnd cell_6t
Xbit_r36_c1 bl_1 br_1 wl_36 vdd gnd cell_6t
Xbit_r37_c1 bl_1 br_1 wl_37 vdd gnd cell_6t
Xbit_r38_c1 bl_1 br_1 wl_38 vdd gnd cell_6t
Xbit_r39_c1 bl_1 br_1 wl_39 vdd gnd cell_6t
Xbit_r40_c1 bl_1 br_1 wl_40 vdd gnd cell_6t
Xbit_r41_c1 bl_1 br_1 wl_41 vdd gnd cell_6t
Xbit_r42_c1 bl_1 br_1 wl_42 vdd gnd cell_6t
Xbit_r43_c1 bl_1 br_1 wl_43 vdd gnd cell_6t
Xbit_r44_c1 bl_1 br_1 wl_44 vdd gnd cell_6t
Xbit_r45_c1 bl_1 br_1 wl_45 vdd gnd cell_6t
Xbit_r46_c1 bl_1 br_1 wl_46 vdd gnd cell_6t
Xbit_r47_c1 bl_1 br_1 wl_47 vdd gnd cell_6t
Xbit_r48_c1 bl_1 br_1 wl_48 vdd gnd cell_6t
Xbit_r49_c1 bl_1 br_1 wl_49 vdd gnd cell_6t
Xbit_r50_c1 bl_1 br_1 wl_50 vdd gnd cell_6t
Xbit_r51_c1 bl_1 br_1 wl_51 vdd gnd cell_6t
Xbit_r52_c1 bl_1 br_1 wl_52 vdd gnd cell_6t
Xbit_r53_c1 bl_1 br_1 wl_53 vdd gnd cell_6t
Xbit_r54_c1 bl_1 br_1 wl_54 vdd gnd cell_6t
Xbit_r55_c1 bl_1 br_1 wl_55 vdd gnd cell_6t
Xbit_r56_c1 bl_1 br_1 wl_56 vdd gnd cell_6t
Xbit_r57_c1 bl_1 br_1 wl_57 vdd gnd cell_6t
Xbit_r58_c1 bl_1 br_1 wl_58 vdd gnd cell_6t
Xbit_r59_c1 bl_1 br_1 wl_59 vdd gnd cell_6t
Xbit_r60_c1 bl_1 br_1 wl_60 vdd gnd cell_6t
Xbit_r61_c1 bl_1 br_1 wl_61 vdd gnd cell_6t
Xbit_r62_c1 bl_1 br_1 wl_62 vdd gnd cell_6t
Xbit_r63_c1 bl_1 br_1 wl_63 vdd gnd cell_6t
Xbit_r64_c1 bl_1 br_1 wl_64 vdd gnd cell_6t
Xbit_r65_c1 bl_1 br_1 wl_65 vdd gnd cell_6t
Xbit_r66_c1 bl_1 br_1 wl_66 vdd gnd cell_6t
Xbit_r67_c1 bl_1 br_1 wl_67 vdd gnd cell_6t
Xbit_r68_c1 bl_1 br_1 wl_68 vdd gnd cell_6t
Xbit_r69_c1 bl_1 br_1 wl_69 vdd gnd cell_6t
Xbit_r70_c1 bl_1 br_1 wl_70 vdd gnd cell_6t
Xbit_r71_c1 bl_1 br_1 wl_71 vdd gnd cell_6t
Xbit_r72_c1 bl_1 br_1 wl_72 vdd gnd cell_6t
Xbit_r73_c1 bl_1 br_1 wl_73 vdd gnd cell_6t
Xbit_r74_c1 bl_1 br_1 wl_74 vdd gnd cell_6t
Xbit_r75_c1 bl_1 br_1 wl_75 vdd gnd cell_6t
Xbit_r76_c1 bl_1 br_1 wl_76 vdd gnd cell_6t
Xbit_r77_c1 bl_1 br_1 wl_77 vdd gnd cell_6t
Xbit_r78_c1 bl_1 br_1 wl_78 vdd gnd cell_6t
Xbit_r79_c1 bl_1 br_1 wl_79 vdd gnd cell_6t
Xbit_r80_c1 bl_1 br_1 wl_80 vdd gnd cell_6t
Xbit_r81_c1 bl_1 br_1 wl_81 vdd gnd cell_6t
Xbit_r82_c1 bl_1 br_1 wl_82 vdd gnd cell_6t
Xbit_r83_c1 bl_1 br_1 wl_83 vdd gnd cell_6t
Xbit_r84_c1 bl_1 br_1 wl_84 vdd gnd cell_6t
Xbit_r85_c1 bl_1 br_1 wl_85 vdd gnd cell_6t
Xbit_r86_c1 bl_1 br_1 wl_86 vdd gnd cell_6t
Xbit_r87_c1 bl_1 br_1 wl_87 vdd gnd cell_6t
Xbit_r88_c1 bl_1 br_1 wl_88 vdd gnd cell_6t
Xbit_r89_c1 bl_1 br_1 wl_89 vdd gnd cell_6t
Xbit_r90_c1 bl_1 br_1 wl_90 vdd gnd cell_6t
Xbit_r91_c1 bl_1 br_1 wl_91 vdd gnd cell_6t
Xbit_r92_c1 bl_1 br_1 wl_92 vdd gnd cell_6t
Xbit_r93_c1 bl_1 br_1 wl_93 vdd gnd cell_6t
Xbit_r94_c1 bl_1 br_1 wl_94 vdd gnd cell_6t
Xbit_r95_c1 bl_1 br_1 wl_95 vdd gnd cell_6t
Xbit_r96_c1 bl_1 br_1 wl_96 vdd gnd cell_6t
Xbit_r97_c1 bl_1 br_1 wl_97 vdd gnd cell_6t
Xbit_r98_c1 bl_1 br_1 wl_98 vdd gnd cell_6t
Xbit_r99_c1 bl_1 br_1 wl_99 vdd gnd cell_6t
Xbit_r100_c1 bl_1 br_1 wl_100 vdd gnd cell_6t
Xbit_r101_c1 bl_1 br_1 wl_101 vdd gnd cell_6t
Xbit_r102_c1 bl_1 br_1 wl_102 vdd gnd cell_6t
Xbit_r103_c1 bl_1 br_1 wl_103 vdd gnd cell_6t
Xbit_r104_c1 bl_1 br_1 wl_104 vdd gnd cell_6t
Xbit_r105_c1 bl_1 br_1 wl_105 vdd gnd cell_6t
Xbit_r106_c1 bl_1 br_1 wl_106 vdd gnd cell_6t
Xbit_r107_c1 bl_1 br_1 wl_107 vdd gnd cell_6t
Xbit_r108_c1 bl_1 br_1 wl_108 vdd gnd cell_6t
Xbit_r109_c1 bl_1 br_1 wl_109 vdd gnd cell_6t
Xbit_r110_c1 bl_1 br_1 wl_110 vdd gnd cell_6t
Xbit_r111_c1 bl_1 br_1 wl_111 vdd gnd cell_6t
Xbit_r112_c1 bl_1 br_1 wl_112 vdd gnd cell_6t
Xbit_r113_c1 bl_1 br_1 wl_113 vdd gnd cell_6t
Xbit_r114_c1 bl_1 br_1 wl_114 vdd gnd cell_6t
Xbit_r115_c1 bl_1 br_1 wl_115 vdd gnd cell_6t
Xbit_r116_c1 bl_1 br_1 wl_116 vdd gnd cell_6t
Xbit_r117_c1 bl_1 br_1 wl_117 vdd gnd cell_6t
Xbit_r118_c1 bl_1 br_1 wl_118 vdd gnd cell_6t
Xbit_r119_c1 bl_1 br_1 wl_119 vdd gnd cell_6t
Xbit_r120_c1 bl_1 br_1 wl_120 vdd gnd cell_6t
Xbit_r121_c1 bl_1 br_1 wl_121 vdd gnd cell_6t
Xbit_r122_c1 bl_1 br_1 wl_122 vdd gnd cell_6t
Xbit_r123_c1 bl_1 br_1 wl_123 vdd gnd cell_6t
Xbit_r124_c1 bl_1 br_1 wl_124 vdd gnd cell_6t
Xbit_r125_c1 bl_1 br_1 wl_125 vdd gnd cell_6t
Xbit_r126_c1 bl_1 br_1 wl_126 vdd gnd cell_6t
Xbit_r127_c1 bl_1 br_1 wl_127 vdd gnd cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd cell_6t
Xbit_r1_c2 bl_2 br_2 wl_1 vdd gnd cell_6t
Xbit_r2_c2 bl_2 br_2 wl_2 vdd gnd cell_6t
Xbit_r3_c2 bl_2 br_2 wl_3 vdd gnd cell_6t
Xbit_r4_c2 bl_2 br_2 wl_4 vdd gnd cell_6t
Xbit_r5_c2 bl_2 br_2 wl_5 vdd gnd cell_6t
Xbit_r6_c2 bl_2 br_2 wl_6 vdd gnd cell_6t
Xbit_r7_c2 bl_2 br_2 wl_7 vdd gnd cell_6t
Xbit_r8_c2 bl_2 br_2 wl_8 vdd gnd cell_6t
Xbit_r9_c2 bl_2 br_2 wl_9 vdd gnd cell_6t
Xbit_r10_c2 bl_2 br_2 wl_10 vdd gnd cell_6t
Xbit_r11_c2 bl_2 br_2 wl_11 vdd gnd cell_6t
Xbit_r12_c2 bl_2 br_2 wl_12 vdd gnd cell_6t
Xbit_r13_c2 bl_2 br_2 wl_13 vdd gnd cell_6t
Xbit_r14_c2 bl_2 br_2 wl_14 vdd gnd cell_6t
Xbit_r15_c2 bl_2 br_2 wl_15 vdd gnd cell_6t
Xbit_r16_c2 bl_2 br_2 wl_16 vdd gnd cell_6t
Xbit_r17_c2 bl_2 br_2 wl_17 vdd gnd cell_6t
Xbit_r18_c2 bl_2 br_2 wl_18 vdd gnd cell_6t
Xbit_r19_c2 bl_2 br_2 wl_19 vdd gnd cell_6t
Xbit_r20_c2 bl_2 br_2 wl_20 vdd gnd cell_6t
Xbit_r21_c2 bl_2 br_2 wl_21 vdd gnd cell_6t
Xbit_r22_c2 bl_2 br_2 wl_22 vdd gnd cell_6t
Xbit_r23_c2 bl_2 br_2 wl_23 vdd gnd cell_6t
Xbit_r24_c2 bl_2 br_2 wl_24 vdd gnd cell_6t
Xbit_r25_c2 bl_2 br_2 wl_25 vdd gnd cell_6t
Xbit_r26_c2 bl_2 br_2 wl_26 vdd gnd cell_6t
Xbit_r27_c2 bl_2 br_2 wl_27 vdd gnd cell_6t
Xbit_r28_c2 bl_2 br_2 wl_28 vdd gnd cell_6t
Xbit_r29_c2 bl_2 br_2 wl_29 vdd gnd cell_6t
Xbit_r30_c2 bl_2 br_2 wl_30 vdd gnd cell_6t
Xbit_r31_c2 bl_2 br_2 wl_31 vdd gnd cell_6t
Xbit_r32_c2 bl_2 br_2 wl_32 vdd gnd cell_6t
Xbit_r33_c2 bl_2 br_2 wl_33 vdd gnd cell_6t
Xbit_r34_c2 bl_2 br_2 wl_34 vdd gnd cell_6t
Xbit_r35_c2 bl_2 br_2 wl_35 vdd gnd cell_6t
Xbit_r36_c2 bl_2 br_2 wl_36 vdd gnd cell_6t
Xbit_r37_c2 bl_2 br_2 wl_37 vdd gnd cell_6t
Xbit_r38_c2 bl_2 br_2 wl_38 vdd gnd cell_6t
Xbit_r39_c2 bl_2 br_2 wl_39 vdd gnd cell_6t
Xbit_r40_c2 bl_2 br_2 wl_40 vdd gnd cell_6t
Xbit_r41_c2 bl_2 br_2 wl_41 vdd gnd cell_6t
Xbit_r42_c2 bl_2 br_2 wl_42 vdd gnd cell_6t
Xbit_r43_c2 bl_2 br_2 wl_43 vdd gnd cell_6t
Xbit_r44_c2 bl_2 br_2 wl_44 vdd gnd cell_6t
Xbit_r45_c2 bl_2 br_2 wl_45 vdd gnd cell_6t
Xbit_r46_c2 bl_2 br_2 wl_46 vdd gnd cell_6t
Xbit_r47_c2 bl_2 br_2 wl_47 vdd gnd cell_6t
Xbit_r48_c2 bl_2 br_2 wl_48 vdd gnd cell_6t
Xbit_r49_c2 bl_2 br_2 wl_49 vdd gnd cell_6t
Xbit_r50_c2 bl_2 br_2 wl_50 vdd gnd cell_6t
Xbit_r51_c2 bl_2 br_2 wl_51 vdd gnd cell_6t
Xbit_r52_c2 bl_2 br_2 wl_52 vdd gnd cell_6t
Xbit_r53_c2 bl_2 br_2 wl_53 vdd gnd cell_6t
Xbit_r54_c2 bl_2 br_2 wl_54 vdd gnd cell_6t
Xbit_r55_c2 bl_2 br_2 wl_55 vdd gnd cell_6t
Xbit_r56_c2 bl_2 br_2 wl_56 vdd gnd cell_6t
Xbit_r57_c2 bl_2 br_2 wl_57 vdd gnd cell_6t
Xbit_r58_c2 bl_2 br_2 wl_58 vdd gnd cell_6t
Xbit_r59_c2 bl_2 br_2 wl_59 vdd gnd cell_6t
Xbit_r60_c2 bl_2 br_2 wl_60 vdd gnd cell_6t
Xbit_r61_c2 bl_2 br_2 wl_61 vdd gnd cell_6t
Xbit_r62_c2 bl_2 br_2 wl_62 vdd gnd cell_6t
Xbit_r63_c2 bl_2 br_2 wl_63 vdd gnd cell_6t
Xbit_r64_c2 bl_2 br_2 wl_64 vdd gnd cell_6t
Xbit_r65_c2 bl_2 br_2 wl_65 vdd gnd cell_6t
Xbit_r66_c2 bl_2 br_2 wl_66 vdd gnd cell_6t
Xbit_r67_c2 bl_2 br_2 wl_67 vdd gnd cell_6t
Xbit_r68_c2 bl_2 br_2 wl_68 vdd gnd cell_6t
Xbit_r69_c2 bl_2 br_2 wl_69 vdd gnd cell_6t
Xbit_r70_c2 bl_2 br_2 wl_70 vdd gnd cell_6t
Xbit_r71_c2 bl_2 br_2 wl_71 vdd gnd cell_6t
Xbit_r72_c2 bl_2 br_2 wl_72 vdd gnd cell_6t
Xbit_r73_c2 bl_2 br_2 wl_73 vdd gnd cell_6t
Xbit_r74_c2 bl_2 br_2 wl_74 vdd gnd cell_6t
Xbit_r75_c2 bl_2 br_2 wl_75 vdd gnd cell_6t
Xbit_r76_c2 bl_2 br_2 wl_76 vdd gnd cell_6t
Xbit_r77_c2 bl_2 br_2 wl_77 vdd gnd cell_6t
Xbit_r78_c2 bl_2 br_2 wl_78 vdd gnd cell_6t
Xbit_r79_c2 bl_2 br_2 wl_79 vdd gnd cell_6t
Xbit_r80_c2 bl_2 br_2 wl_80 vdd gnd cell_6t
Xbit_r81_c2 bl_2 br_2 wl_81 vdd gnd cell_6t
Xbit_r82_c2 bl_2 br_2 wl_82 vdd gnd cell_6t
Xbit_r83_c2 bl_2 br_2 wl_83 vdd gnd cell_6t
Xbit_r84_c2 bl_2 br_2 wl_84 vdd gnd cell_6t
Xbit_r85_c2 bl_2 br_2 wl_85 vdd gnd cell_6t
Xbit_r86_c2 bl_2 br_2 wl_86 vdd gnd cell_6t
Xbit_r87_c2 bl_2 br_2 wl_87 vdd gnd cell_6t
Xbit_r88_c2 bl_2 br_2 wl_88 vdd gnd cell_6t
Xbit_r89_c2 bl_2 br_2 wl_89 vdd gnd cell_6t
Xbit_r90_c2 bl_2 br_2 wl_90 vdd gnd cell_6t
Xbit_r91_c2 bl_2 br_2 wl_91 vdd gnd cell_6t
Xbit_r92_c2 bl_2 br_2 wl_92 vdd gnd cell_6t
Xbit_r93_c2 bl_2 br_2 wl_93 vdd gnd cell_6t
Xbit_r94_c2 bl_2 br_2 wl_94 vdd gnd cell_6t
Xbit_r95_c2 bl_2 br_2 wl_95 vdd gnd cell_6t
Xbit_r96_c2 bl_2 br_2 wl_96 vdd gnd cell_6t
Xbit_r97_c2 bl_2 br_2 wl_97 vdd gnd cell_6t
Xbit_r98_c2 bl_2 br_2 wl_98 vdd gnd cell_6t
Xbit_r99_c2 bl_2 br_2 wl_99 vdd gnd cell_6t
Xbit_r100_c2 bl_2 br_2 wl_100 vdd gnd cell_6t
Xbit_r101_c2 bl_2 br_2 wl_101 vdd gnd cell_6t
Xbit_r102_c2 bl_2 br_2 wl_102 vdd gnd cell_6t
Xbit_r103_c2 bl_2 br_2 wl_103 vdd gnd cell_6t
Xbit_r104_c2 bl_2 br_2 wl_104 vdd gnd cell_6t
Xbit_r105_c2 bl_2 br_2 wl_105 vdd gnd cell_6t
Xbit_r106_c2 bl_2 br_2 wl_106 vdd gnd cell_6t
Xbit_r107_c2 bl_2 br_2 wl_107 vdd gnd cell_6t
Xbit_r108_c2 bl_2 br_2 wl_108 vdd gnd cell_6t
Xbit_r109_c2 bl_2 br_2 wl_109 vdd gnd cell_6t
Xbit_r110_c2 bl_2 br_2 wl_110 vdd gnd cell_6t
Xbit_r111_c2 bl_2 br_2 wl_111 vdd gnd cell_6t
Xbit_r112_c2 bl_2 br_2 wl_112 vdd gnd cell_6t
Xbit_r113_c2 bl_2 br_2 wl_113 vdd gnd cell_6t
Xbit_r114_c2 bl_2 br_2 wl_114 vdd gnd cell_6t
Xbit_r115_c2 bl_2 br_2 wl_115 vdd gnd cell_6t
Xbit_r116_c2 bl_2 br_2 wl_116 vdd gnd cell_6t
Xbit_r117_c2 bl_2 br_2 wl_117 vdd gnd cell_6t
Xbit_r118_c2 bl_2 br_2 wl_118 vdd gnd cell_6t
Xbit_r119_c2 bl_2 br_2 wl_119 vdd gnd cell_6t
Xbit_r120_c2 bl_2 br_2 wl_120 vdd gnd cell_6t
Xbit_r121_c2 bl_2 br_2 wl_121 vdd gnd cell_6t
Xbit_r122_c2 bl_2 br_2 wl_122 vdd gnd cell_6t
Xbit_r123_c2 bl_2 br_2 wl_123 vdd gnd cell_6t
Xbit_r124_c2 bl_2 br_2 wl_124 vdd gnd cell_6t
Xbit_r125_c2 bl_2 br_2 wl_125 vdd gnd cell_6t
Xbit_r126_c2 bl_2 br_2 wl_126 vdd gnd cell_6t
Xbit_r127_c2 bl_2 br_2 wl_127 vdd gnd cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd cell_6t
Xbit_r1_c3 bl_3 br_3 wl_1 vdd gnd cell_6t
Xbit_r2_c3 bl_3 br_3 wl_2 vdd gnd cell_6t
Xbit_r3_c3 bl_3 br_3 wl_3 vdd gnd cell_6t
Xbit_r4_c3 bl_3 br_3 wl_4 vdd gnd cell_6t
Xbit_r5_c3 bl_3 br_3 wl_5 vdd gnd cell_6t
Xbit_r6_c3 bl_3 br_3 wl_6 vdd gnd cell_6t
Xbit_r7_c3 bl_3 br_3 wl_7 vdd gnd cell_6t
Xbit_r8_c3 bl_3 br_3 wl_8 vdd gnd cell_6t
Xbit_r9_c3 bl_3 br_3 wl_9 vdd gnd cell_6t
Xbit_r10_c3 bl_3 br_3 wl_10 vdd gnd cell_6t
Xbit_r11_c3 bl_3 br_3 wl_11 vdd gnd cell_6t
Xbit_r12_c3 bl_3 br_3 wl_12 vdd gnd cell_6t
Xbit_r13_c3 bl_3 br_3 wl_13 vdd gnd cell_6t
Xbit_r14_c3 bl_3 br_3 wl_14 vdd gnd cell_6t
Xbit_r15_c3 bl_3 br_3 wl_15 vdd gnd cell_6t
Xbit_r16_c3 bl_3 br_3 wl_16 vdd gnd cell_6t
Xbit_r17_c3 bl_3 br_3 wl_17 vdd gnd cell_6t
Xbit_r18_c3 bl_3 br_3 wl_18 vdd gnd cell_6t
Xbit_r19_c3 bl_3 br_3 wl_19 vdd gnd cell_6t
Xbit_r20_c3 bl_3 br_3 wl_20 vdd gnd cell_6t
Xbit_r21_c3 bl_3 br_3 wl_21 vdd gnd cell_6t
Xbit_r22_c3 bl_3 br_3 wl_22 vdd gnd cell_6t
Xbit_r23_c3 bl_3 br_3 wl_23 vdd gnd cell_6t
Xbit_r24_c3 bl_3 br_3 wl_24 vdd gnd cell_6t
Xbit_r25_c3 bl_3 br_3 wl_25 vdd gnd cell_6t
Xbit_r26_c3 bl_3 br_3 wl_26 vdd gnd cell_6t
Xbit_r27_c3 bl_3 br_3 wl_27 vdd gnd cell_6t
Xbit_r28_c3 bl_3 br_3 wl_28 vdd gnd cell_6t
Xbit_r29_c3 bl_3 br_3 wl_29 vdd gnd cell_6t
Xbit_r30_c3 bl_3 br_3 wl_30 vdd gnd cell_6t
Xbit_r31_c3 bl_3 br_3 wl_31 vdd gnd cell_6t
Xbit_r32_c3 bl_3 br_3 wl_32 vdd gnd cell_6t
Xbit_r33_c3 bl_3 br_3 wl_33 vdd gnd cell_6t
Xbit_r34_c3 bl_3 br_3 wl_34 vdd gnd cell_6t
Xbit_r35_c3 bl_3 br_3 wl_35 vdd gnd cell_6t
Xbit_r36_c3 bl_3 br_3 wl_36 vdd gnd cell_6t
Xbit_r37_c3 bl_3 br_3 wl_37 vdd gnd cell_6t
Xbit_r38_c3 bl_3 br_3 wl_38 vdd gnd cell_6t
Xbit_r39_c3 bl_3 br_3 wl_39 vdd gnd cell_6t
Xbit_r40_c3 bl_3 br_3 wl_40 vdd gnd cell_6t
Xbit_r41_c3 bl_3 br_3 wl_41 vdd gnd cell_6t
Xbit_r42_c3 bl_3 br_3 wl_42 vdd gnd cell_6t
Xbit_r43_c3 bl_3 br_3 wl_43 vdd gnd cell_6t
Xbit_r44_c3 bl_3 br_3 wl_44 vdd gnd cell_6t
Xbit_r45_c3 bl_3 br_3 wl_45 vdd gnd cell_6t
Xbit_r46_c3 bl_3 br_3 wl_46 vdd gnd cell_6t
Xbit_r47_c3 bl_3 br_3 wl_47 vdd gnd cell_6t
Xbit_r48_c3 bl_3 br_3 wl_48 vdd gnd cell_6t
Xbit_r49_c3 bl_3 br_3 wl_49 vdd gnd cell_6t
Xbit_r50_c3 bl_3 br_3 wl_50 vdd gnd cell_6t
Xbit_r51_c3 bl_3 br_3 wl_51 vdd gnd cell_6t
Xbit_r52_c3 bl_3 br_3 wl_52 vdd gnd cell_6t
Xbit_r53_c3 bl_3 br_3 wl_53 vdd gnd cell_6t
Xbit_r54_c3 bl_3 br_3 wl_54 vdd gnd cell_6t
Xbit_r55_c3 bl_3 br_3 wl_55 vdd gnd cell_6t
Xbit_r56_c3 bl_3 br_3 wl_56 vdd gnd cell_6t
Xbit_r57_c3 bl_3 br_3 wl_57 vdd gnd cell_6t
Xbit_r58_c3 bl_3 br_3 wl_58 vdd gnd cell_6t
Xbit_r59_c3 bl_3 br_3 wl_59 vdd gnd cell_6t
Xbit_r60_c3 bl_3 br_3 wl_60 vdd gnd cell_6t
Xbit_r61_c3 bl_3 br_3 wl_61 vdd gnd cell_6t
Xbit_r62_c3 bl_3 br_3 wl_62 vdd gnd cell_6t
Xbit_r63_c3 bl_3 br_3 wl_63 vdd gnd cell_6t
Xbit_r64_c3 bl_3 br_3 wl_64 vdd gnd cell_6t
Xbit_r65_c3 bl_3 br_3 wl_65 vdd gnd cell_6t
Xbit_r66_c3 bl_3 br_3 wl_66 vdd gnd cell_6t
Xbit_r67_c3 bl_3 br_3 wl_67 vdd gnd cell_6t
Xbit_r68_c3 bl_3 br_3 wl_68 vdd gnd cell_6t
Xbit_r69_c3 bl_3 br_3 wl_69 vdd gnd cell_6t
Xbit_r70_c3 bl_3 br_3 wl_70 vdd gnd cell_6t
Xbit_r71_c3 bl_3 br_3 wl_71 vdd gnd cell_6t
Xbit_r72_c3 bl_3 br_3 wl_72 vdd gnd cell_6t
Xbit_r73_c3 bl_3 br_3 wl_73 vdd gnd cell_6t
Xbit_r74_c3 bl_3 br_3 wl_74 vdd gnd cell_6t
Xbit_r75_c3 bl_3 br_3 wl_75 vdd gnd cell_6t
Xbit_r76_c3 bl_3 br_3 wl_76 vdd gnd cell_6t
Xbit_r77_c3 bl_3 br_3 wl_77 vdd gnd cell_6t
Xbit_r78_c3 bl_3 br_3 wl_78 vdd gnd cell_6t
Xbit_r79_c3 bl_3 br_3 wl_79 vdd gnd cell_6t
Xbit_r80_c3 bl_3 br_3 wl_80 vdd gnd cell_6t
Xbit_r81_c3 bl_3 br_3 wl_81 vdd gnd cell_6t
Xbit_r82_c3 bl_3 br_3 wl_82 vdd gnd cell_6t
Xbit_r83_c3 bl_3 br_3 wl_83 vdd gnd cell_6t
Xbit_r84_c3 bl_3 br_3 wl_84 vdd gnd cell_6t
Xbit_r85_c3 bl_3 br_3 wl_85 vdd gnd cell_6t
Xbit_r86_c3 bl_3 br_3 wl_86 vdd gnd cell_6t
Xbit_r87_c3 bl_3 br_3 wl_87 vdd gnd cell_6t
Xbit_r88_c3 bl_3 br_3 wl_88 vdd gnd cell_6t
Xbit_r89_c3 bl_3 br_3 wl_89 vdd gnd cell_6t
Xbit_r90_c3 bl_3 br_3 wl_90 vdd gnd cell_6t
Xbit_r91_c3 bl_3 br_3 wl_91 vdd gnd cell_6t
Xbit_r92_c3 bl_3 br_3 wl_92 vdd gnd cell_6t
Xbit_r93_c3 bl_3 br_3 wl_93 vdd gnd cell_6t
Xbit_r94_c3 bl_3 br_3 wl_94 vdd gnd cell_6t
Xbit_r95_c3 bl_3 br_3 wl_95 vdd gnd cell_6t
Xbit_r96_c3 bl_3 br_3 wl_96 vdd gnd cell_6t
Xbit_r97_c3 bl_3 br_3 wl_97 vdd gnd cell_6t
Xbit_r98_c3 bl_3 br_3 wl_98 vdd gnd cell_6t
Xbit_r99_c3 bl_3 br_3 wl_99 vdd gnd cell_6t
Xbit_r100_c3 bl_3 br_3 wl_100 vdd gnd cell_6t
Xbit_r101_c3 bl_3 br_3 wl_101 vdd gnd cell_6t
Xbit_r102_c3 bl_3 br_3 wl_102 vdd gnd cell_6t
Xbit_r103_c3 bl_3 br_3 wl_103 vdd gnd cell_6t
Xbit_r104_c3 bl_3 br_3 wl_104 vdd gnd cell_6t
Xbit_r105_c3 bl_3 br_3 wl_105 vdd gnd cell_6t
Xbit_r106_c3 bl_3 br_3 wl_106 vdd gnd cell_6t
Xbit_r107_c3 bl_3 br_3 wl_107 vdd gnd cell_6t
Xbit_r108_c3 bl_3 br_3 wl_108 vdd gnd cell_6t
Xbit_r109_c3 bl_3 br_3 wl_109 vdd gnd cell_6t
Xbit_r110_c3 bl_3 br_3 wl_110 vdd gnd cell_6t
Xbit_r111_c3 bl_3 br_3 wl_111 vdd gnd cell_6t
Xbit_r112_c3 bl_3 br_3 wl_112 vdd gnd cell_6t
Xbit_r113_c3 bl_3 br_3 wl_113 vdd gnd cell_6t
Xbit_r114_c3 bl_3 br_3 wl_114 vdd gnd cell_6t
Xbit_r115_c3 bl_3 br_3 wl_115 vdd gnd cell_6t
Xbit_r116_c3 bl_3 br_3 wl_116 vdd gnd cell_6t
Xbit_r117_c3 bl_3 br_3 wl_117 vdd gnd cell_6t
Xbit_r118_c3 bl_3 br_3 wl_118 vdd gnd cell_6t
Xbit_r119_c3 bl_3 br_3 wl_119 vdd gnd cell_6t
Xbit_r120_c3 bl_3 br_3 wl_120 vdd gnd cell_6t
Xbit_r121_c3 bl_3 br_3 wl_121 vdd gnd cell_6t
Xbit_r122_c3 bl_3 br_3 wl_122 vdd gnd cell_6t
Xbit_r123_c3 bl_3 br_3 wl_123 vdd gnd cell_6t
Xbit_r124_c3 bl_3 br_3 wl_124 vdd gnd cell_6t
Xbit_r125_c3 bl_3 br_3 wl_125 vdd gnd cell_6t
Xbit_r126_c3 bl_3 br_3 wl_126 vdd gnd cell_6t
Xbit_r127_c3 bl_3 br_3 wl_127 vdd gnd cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd cell_6t
Xbit_r1_c4 bl_4 br_4 wl_1 vdd gnd cell_6t
Xbit_r2_c4 bl_4 br_4 wl_2 vdd gnd cell_6t
Xbit_r3_c4 bl_4 br_4 wl_3 vdd gnd cell_6t
Xbit_r4_c4 bl_4 br_4 wl_4 vdd gnd cell_6t
Xbit_r5_c4 bl_4 br_4 wl_5 vdd gnd cell_6t
Xbit_r6_c4 bl_4 br_4 wl_6 vdd gnd cell_6t
Xbit_r7_c4 bl_4 br_4 wl_7 vdd gnd cell_6t
Xbit_r8_c4 bl_4 br_4 wl_8 vdd gnd cell_6t
Xbit_r9_c4 bl_4 br_4 wl_9 vdd gnd cell_6t
Xbit_r10_c4 bl_4 br_4 wl_10 vdd gnd cell_6t
Xbit_r11_c4 bl_4 br_4 wl_11 vdd gnd cell_6t
Xbit_r12_c4 bl_4 br_4 wl_12 vdd gnd cell_6t
Xbit_r13_c4 bl_4 br_4 wl_13 vdd gnd cell_6t
Xbit_r14_c4 bl_4 br_4 wl_14 vdd gnd cell_6t
Xbit_r15_c4 bl_4 br_4 wl_15 vdd gnd cell_6t
Xbit_r16_c4 bl_4 br_4 wl_16 vdd gnd cell_6t
Xbit_r17_c4 bl_4 br_4 wl_17 vdd gnd cell_6t
Xbit_r18_c4 bl_4 br_4 wl_18 vdd gnd cell_6t
Xbit_r19_c4 bl_4 br_4 wl_19 vdd gnd cell_6t
Xbit_r20_c4 bl_4 br_4 wl_20 vdd gnd cell_6t
Xbit_r21_c4 bl_4 br_4 wl_21 vdd gnd cell_6t
Xbit_r22_c4 bl_4 br_4 wl_22 vdd gnd cell_6t
Xbit_r23_c4 bl_4 br_4 wl_23 vdd gnd cell_6t
Xbit_r24_c4 bl_4 br_4 wl_24 vdd gnd cell_6t
Xbit_r25_c4 bl_4 br_4 wl_25 vdd gnd cell_6t
Xbit_r26_c4 bl_4 br_4 wl_26 vdd gnd cell_6t
Xbit_r27_c4 bl_4 br_4 wl_27 vdd gnd cell_6t
Xbit_r28_c4 bl_4 br_4 wl_28 vdd gnd cell_6t
Xbit_r29_c4 bl_4 br_4 wl_29 vdd gnd cell_6t
Xbit_r30_c4 bl_4 br_4 wl_30 vdd gnd cell_6t
Xbit_r31_c4 bl_4 br_4 wl_31 vdd gnd cell_6t
Xbit_r32_c4 bl_4 br_4 wl_32 vdd gnd cell_6t
Xbit_r33_c4 bl_4 br_4 wl_33 vdd gnd cell_6t
Xbit_r34_c4 bl_4 br_4 wl_34 vdd gnd cell_6t
Xbit_r35_c4 bl_4 br_4 wl_35 vdd gnd cell_6t
Xbit_r36_c4 bl_4 br_4 wl_36 vdd gnd cell_6t
Xbit_r37_c4 bl_4 br_4 wl_37 vdd gnd cell_6t
Xbit_r38_c4 bl_4 br_4 wl_38 vdd gnd cell_6t
Xbit_r39_c4 bl_4 br_4 wl_39 vdd gnd cell_6t
Xbit_r40_c4 bl_4 br_4 wl_40 vdd gnd cell_6t
Xbit_r41_c4 bl_4 br_4 wl_41 vdd gnd cell_6t
Xbit_r42_c4 bl_4 br_4 wl_42 vdd gnd cell_6t
Xbit_r43_c4 bl_4 br_4 wl_43 vdd gnd cell_6t
Xbit_r44_c4 bl_4 br_4 wl_44 vdd gnd cell_6t
Xbit_r45_c4 bl_4 br_4 wl_45 vdd gnd cell_6t
Xbit_r46_c4 bl_4 br_4 wl_46 vdd gnd cell_6t
Xbit_r47_c4 bl_4 br_4 wl_47 vdd gnd cell_6t
Xbit_r48_c4 bl_4 br_4 wl_48 vdd gnd cell_6t
Xbit_r49_c4 bl_4 br_4 wl_49 vdd gnd cell_6t
Xbit_r50_c4 bl_4 br_4 wl_50 vdd gnd cell_6t
Xbit_r51_c4 bl_4 br_4 wl_51 vdd gnd cell_6t
Xbit_r52_c4 bl_4 br_4 wl_52 vdd gnd cell_6t
Xbit_r53_c4 bl_4 br_4 wl_53 vdd gnd cell_6t
Xbit_r54_c4 bl_4 br_4 wl_54 vdd gnd cell_6t
Xbit_r55_c4 bl_4 br_4 wl_55 vdd gnd cell_6t
Xbit_r56_c4 bl_4 br_4 wl_56 vdd gnd cell_6t
Xbit_r57_c4 bl_4 br_4 wl_57 vdd gnd cell_6t
Xbit_r58_c4 bl_4 br_4 wl_58 vdd gnd cell_6t
Xbit_r59_c4 bl_4 br_4 wl_59 vdd gnd cell_6t
Xbit_r60_c4 bl_4 br_4 wl_60 vdd gnd cell_6t
Xbit_r61_c4 bl_4 br_4 wl_61 vdd gnd cell_6t
Xbit_r62_c4 bl_4 br_4 wl_62 vdd gnd cell_6t
Xbit_r63_c4 bl_4 br_4 wl_63 vdd gnd cell_6t
Xbit_r64_c4 bl_4 br_4 wl_64 vdd gnd cell_6t
Xbit_r65_c4 bl_4 br_4 wl_65 vdd gnd cell_6t
Xbit_r66_c4 bl_4 br_4 wl_66 vdd gnd cell_6t
Xbit_r67_c4 bl_4 br_4 wl_67 vdd gnd cell_6t
Xbit_r68_c4 bl_4 br_4 wl_68 vdd gnd cell_6t
Xbit_r69_c4 bl_4 br_4 wl_69 vdd gnd cell_6t
Xbit_r70_c4 bl_4 br_4 wl_70 vdd gnd cell_6t
Xbit_r71_c4 bl_4 br_4 wl_71 vdd gnd cell_6t
Xbit_r72_c4 bl_4 br_4 wl_72 vdd gnd cell_6t
Xbit_r73_c4 bl_4 br_4 wl_73 vdd gnd cell_6t
Xbit_r74_c4 bl_4 br_4 wl_74 vdd gnd cell_6t
Xbit_r75_c4 bl_4 br_4 wl_75 vdd gnd cell_6t
Xbit_r76_c4 bl_4 br_4 wl_76 vdd gnd cell_6t
Xbit_r77_c4 bl_4 br_4 wl_77 vdd gnd cell_6t
Xbit_r78_c4 bl_4 br_4 wl_78 vdd gnd cell_6t
Xbit_r79_c4 bl_4 br_4 wl_79 vdd gnd cell_6t
Xbit_r80_c4 bl_4 br_4 wl_80 vdd gnd cell_6t
Xbit_r81_c4 bl_4 br_4 wl_81 vdd gnd cell_6t
Xbit_r82_c4 bl_4 br_4 wl_82 vdd gnd cell_6t
Xbit_r83_c4 bl_4 br_4 wl_83 vdd gnd cell_6t
Xbit_r84_c4 bl_4 br_4 wl_84 vdd gnd cell_6t
Xbit_r85_c4 bl_4 br_4 wl_85 vdd gnd cell_6t
Xbit_r86_c4 bl_4 br_4 wl_86 vdd gnd cell_6t
Xbit_r87_c4 bl_4 br_4 wl_87 vdd gnd cell_6t
Xbit_r88_c4 bl_4 br_4 wl_88 vdd gnd cell_6t
Xbit_r89_c4 bl_4 br_4 wl_89 vdd gnd cell_6t
Xbit_r90_c4 bl_4 br_4 wl_90 vdd gnd cell_6t
Xbit_r91_c4 bl_4 br_4 wl_91 vdd gnd cell_6t
Xbit_r92_c4 bl_4 br_4 wl_92 vdd gnd cell_6t
Xbit_r93_c4 bl_4 br_4 wl_93 vdd gnd cell_6t
Xbit_r94_c4 bl_4 br_4 wl_94 vdd gnd cell_6t
Xbit_r95_c4 bl_4 br_4 wl_95 vdd gnd cell_6t
Xbit_r96_c4 bl_4 br_4 wl_96 vdd gnd cell_6t
Xbit_r97_c4 bl_4 br_4 wl_97 vdd gnd cell_6t
Xbit_r98_c4 bl_4 br_4 wl_98 vdd gnd cell_6t
Xbit_r99_c4 bl_4 br_4 wl_99 vdd gnd cell_6t
Xbit_r100_c4 bl_4 br_4 wl_100 vdd gnd cell_6t
Xbit_r101_c4 bl_4 br_4 wl_101 vdd gnd cell_6t
Xbit_r102_c4 bl_4 br_4 wl_102 vdd gnd cell_6t
Xbit_r103_c4 bl_4 br_4 wl_103 vdd gnd cell_6t
Xbit_r104_c4 bl_4 br_4 wl_104 vdd gnd cell_6t
Xbit_r105_c4 bl_4 br_4 wl_105 vdd gnd cell_6t
Xbit_r106_c4 bl_4 br_4 wl_106 vdd gnd cell_6t
Xbit_r107_c4 bl_4 br_4 wl_107 vdd gnd cell_6t
Xbit_r108_c4 bl_4 br_4 wl_108 vdd gnd cell_6t
Xbit_r109_c4 bl_4 br_4 wl_109 vdd gnd cell_6t
Xbit_r110_c4 bl_4 br_4 wl_110 vdd gnd cell_6t
Xbit_r111_c4 bl_4 br_4 wl_111 vdd gnd cell_6t
Xbit_r112_c4 bl_4 br_4 wl_112 vdd gnd cell_6t
Xbit_r113_c4 bl_4 br_4 wl_113 vdd gnd cell_6t
Xbit_r114_c4 bl_4 br_4 wl_114 vdd gnd cell_6t
Xbit_r115_c4 bl_4 br_4 wl_115 vdd gnd cell_6t
Xbit_r116_c4 bl_4 br_4 wl_116 vdd gnd cell_6t
Xbit_r117_c4 bl_4 br_4 wl_117 vdd gnd cell_6t
Xbit_r118_c4 bl_4 br_4 wl_118 vdd gnd cell_6t
Xbit_r119_c4 bl_4 br_4 wl_119 vdd gnd cell_6t
Xbit_r120_c4 bl_4 br_4 wl_120 vdd gnd cell_6t
Xbit_r121_c4 bl_4 br_4 wl_121 vdd gnd cell_6t
Xbit_r122_c4 bl_4 br_4 wl_122 vdd gnd cell_6t
Xbit_r123_c4 bl_4 br_4 wl_123 vdd gnd cell_6t
Xbit_r124_c4 bl_4 br_4 wl_124 vdd gnd cell_6t
Xbit_r125_c4 bl_4 br_4 wl_125 vdd gnd cell_6t
Xbit_r126_c4 bl_4 br_4 wl_126 vdd gnd cell_6t
Xbit_r127_c4 bl_4 br_4 wl_127 vdd gnd cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd cell_6t
Xbit_r1_c5 bl_5 br_5 wl_1 vdd gnd cell_6t
Xbit_r2_c5 bl_5 br_5 wl_2 vdd gnd cell_6t
Xbit_r3_c5 bl_5 br_5 wl_3 vdd gnd cell_6t
Xbit_r4_c5 bl_5 br_5 wl_4 vdd gnd cell_6t
Xbit_r5_c5 bl_5 br_5 wl_5 vdd gnd cell_6t
Xbit_r6_c5 bl_5 br_5 wl_6 vdd gnd cell_6t
Xbit_r7_c5 bl_5 br_5 wl_7 vdd gnd cell_6t
Xbit_r8_c5 bl_5 br_5 wl_8 vdd gnd cell_6t
Xbit_r9_c5 bl_5 br_5 wl_9 vdd gnd cell_6t
Xbit_r10_c5 bl_5 br_5 wl_10 vdd gnd cell_6t
Xbit_r11_c5 bl_5 br_5 wl_11 vdd gnd cell_6t
Xbit_r12_c5 bl_5 br_5 wl_12 vdd gnd cell_6t
Xbit_r13_c5 bl_5 br_5 wl_13 vdd gnd cell_6t
Xbit_r14_c5 bl_5 br_5 wl_14 vdd gnd cell_6t
Xbit_r15_c5 bl_5 br_5 wl_15 vdd gnd cell_6t
Xbit_r16_c5 bl_5 br_5 wl_16 vdd gnd cell_6t
Xbit_r17_c5 bl_5 br_5 wl_17 vdd gnd cell_6t
Xbit_r18_c5 bl_5 br_5 wl_18 vdd gnd cell_6t
Xbit_r19_c5 bl_5 br_5 wl_19 vdd gnd cell_6t
Xbit_r20_c5 bl_5 br_5 wl_20 vdd gnd cell_6t
Xbit_r21_c5 bl_5 br_5 wl_21 vdd gnd cell_6t
Xbit_r22_c5 bl_5 br_5 wl_22 vdd gnd cell_6t
Xbit_r23_c5 bl_5 br_5 wl_23 vdd gnd cell_6t
Xbit_r24_c5 bl_5 br_5 wl_24 vdd gnd cell_6t
Xbit_r25_c5 bl_5 br_5 wl_25 vdd gnd cell_6t
Xbit_r26_c5 bl_5 br_5 wl_26 vdd gnd cell_6t
Xbit_r27_c5 bl_5 br_5 wl_27 vdd gnd cell_6t
Xbit_r28_c5 bl_5 br_5 wl_28 vdd gnd cell_6t
Xbit_r29_c5 bl_5 br_5 wl_29 vdd gnd cell_6t
Xbit_r30_c5 bl_5 br_5 wl_30 vdd gnd cell_6t
Xbit_r31_c5 bl_5 br_5 wl_31 vdd gnd cell_6t
Xbit_r32_c5 bl_5 br_5 wl_32 vdd gnd cell_6t
Xbit_r33_c5 bl_5 br_5 wl_33 vdd gnd cell_6t
Xbit_r34_c5 bl_5 br_5 wl_34 vdd gnd cell_6t
Xbit_r35_c5 bl_5 br_5 wl_35 vdd gnd cell_6t
Xbit_r36_c5 bl_5 br_5 wl_36 vdd gnd cell_6t
Xbit_r37_c5 bl_5 br_5 wl_37 vdd gnd cell_6t
Xbit_r38_c5 bl_5 br_5 wl_38 vdd gnd cell_6t
Xbit_r39_c5 bl_5 br_5 wl_39 vdd gnd cell_6t
Xbit_r40_c5 bl_5 br_5 wl_40 vdd gnd cell_6t
Xbit_r41_c5 bl_5 br_5 wl_41 vdd gnd cell_6t
Xbit_r42_c5 bl_5 br_5 wl_42 vdd gnd cell_6t
Xbit_r43_c5 bl_5 br_5 wl_43 vdd gnd cell_6t
Xbit_r44_c5 bl_5 br_5 wl_44 vdd gnd cell_6t
Xbit_r45_c5 bl_5 br_5 wl_45 vdd gnd cell_6t
Xbit_r46_c5 bl_5 br_5 wl_46 vdd gnd cell_6t
Xbit_r47_c5 bl_5 br_5 wl_47 vdd gnd cell_6t
Xbit_r48_c5 bl_5 br_5 wl_48 vdd gnd cell_6t
Xbit_r49_c5 bl_5 br_5 wl_49 vdd gnd cell_6t
Xbit_r50_c5 bl_5 br_5 wl_50 vdd gnd cell_6t
Xbit_r51_c5 bl_5 br_5 wl_51 vdd gnd cell_6t
Xbit_r52_c5 bl_5 br_5 wl_52 vdd gnd cell_6t
Xbit_r53_c5 bl_5 br_5 wl_53 vdd gnd cell_6t
Xbit_r54_c5 bl_5 br_5 wl_54 vdd gnd cell_6t
Xbit_r55_c5 bl_5 br_5 wl_55 vdd gnd cell_6t
Xbit_r56_c5 bl_5 br_5 wl_56 vdd gnd cell_6t
Xbit_r57_c5 bl_5 br_5 wl_57 vdd gnd cell_6t
Xbit_r58_c5 bl_5 br_5 wl_58 vdd gnd cell_6t
Xbit_r59_c5 bl_5 br_5 wl_59 vdd gnd cell_6t
Xbit_r60_c5 bl_5 br_5 wl_60 vdd gnd cell_6t
Xbit_r61_c5 bl_5 br_5 wl_61 vdd gnd cell_6t
Xbit_r62_c5 bl_5 br_5 wl_62 vdd gnd cell_6t
Xbit_r63_c5 bl_5 br_5 wl_63 vdd gnd cell_6t
Xbit_r64_c5 bl_5 br_5 wl_64 vdd gnd cell_6t
Xbit_r65_c5 bl_5 br_5 wl_65 vdd gnd cell_6t
Xbit_r66_c5 bl_5 br_5 wl_66 vdd gnd cell_6t
Xbit_r67_c5 bl_5 br_5 wl_67 vdd gnd cell_6t
Xbit_r68_c5 bl_5 br_5 wl_68 vdd gnd cell_6t
Xbit_r69_c5 bl_5 br_5 wl_69 vdd gnd cell_6t
Xbit_r70_c5 bl_5 br_5 wl_70 vdd gnd cell_6t
Xbit_r71_c5 bl_5 br_5 wl_71 vdd gnd cell_6t
Xbit_r72_c5 bl_5 br_5 wl_72 vdd gnd cell_6t
Xbit_r73_c5 bl_5 br_5 wl_73 vdd gnd cell_6t
Xbit_r74_c5 bl_5 br_5 wl_74 vdd gnd cell_6t
Xbit_r75_c5 bl_5 br_5 wl_75 vdd gnd cell_6t
Xbit_r76_c5 bl_5 br_5 wl_76 vdd gnd cell_6t
Xbit_r77_c5 bl_5 br_5 wl_77 vdd gnd cell_6t
Xbit_r78_c5 bl_5 br_5 wl_78 vdd gnd cell_6t
Xbit_r79_c5 bl_5 br_5 wl_79 vdd gnd cell_6t
Xbit_r80_c5 bl_5 br_5 wl_80 vdd gnd cell_6t
Xbit_r81_c5 bl_5 br_5 wl_81 vdd gnd cell_6t
Xbit_r82_c5 bl_5 br_5 wl_82 vdd gnd cell_6t
Xbit_r83_c5 bl_5 br_5 wl_83 vdd gnd cell_6t
Xbit_r84_c5 bl_5 br_5 wl_84 vdd gnd cell_6t
Xbit_r85_c5 bl_5 br_5 wl_85 vdd gnd cell_6t
Xbit_r86_c5 bl_5 br_5 wl_86 vdd gnd cell_6t
Xbit_r87_c5 bl_5 br_5 wl_87 vdd gnd cell_6t
Xbit_r88_c5 bl_5 br_5 wl_88 vdd gnd cell_6t
Xbit_r89_c5 bl_5 br_5 wl_89 vdd gnd cell_6t
Xbit_r90_c5 bl_5 br_5 wl_90 vdd gnd cell_6t
Xbit_r91_c5 bl_5 br_5 wl_91 vdd gnd cell_6t
Xbit_r92_c5 bl_5 br_5 wl_92 vdd gnd cell_6t
Xbit_r93_c5 bl_5 br_5 wl_93 vdd gnd cell_6t
Xbit_r94_c5 bl_5 br_5 wl_94 vdd gnd cell_6t
Xbit_r95_c5 bl_5 br_5 wl_95 vdd gnd cell_6t
Xbit_r96_c5 bl_5 br_5 wl_96 vdd gnd cell_6t
Xbit_r97_c5 bl_5 br_5 wl_97 vdd gnd cell_6t
Xbit_r98_c5 bl_5 br_5 wl_98 vdd gnd cell_6t
Xbit_r99_c5 bl_5 br_5 wl_99 vdd gnd cell_6t
Xbit_r100_c5 bl_5 br_5 wl_100 vdd gnd cell_6t
Xbit_r101_c5 bl_5 br_5 wl_101 vdd gnd cell_6t
Xbit_r102_c5 bl_5 br_5 wl_102 vdd gnd cell_6t
Xbit_r103_c5 bl_5 br_5 wl_103 vdd gnd cell_6t
Xbit_r104_c5 bl_5 br_5 wl_104 vdd gnd cell_6t
Xbit_r105_c5 bl_5 br_5 wl_105 vdd gnd cell_6t
Xbit_r106_c5 bl_5 br_5 wl_106 vdd gnd cell_6t
Xbit_r107_c5 bl_5 br_5 wl_107 vdd gnd cell_6t
Xbit_r108_c5 bl_5 br_5 wl_108 vdd gnd cell_6t
Xbit_r109_c5 bl_5 br_5 wl_109 vdd gnd cell_6t
Xbit_r110_c5 bl_5 br_5 wl_110 vdd gnd cell_6t
Xbit_r111_c5 bl_5 br_5 wl_111 vdd gnd cell_6t
Xbit_r112_c5 bl_5 br_5 wl_112 vdd gnd cell_6t
Xbit_r113_c5 bl_5 br_5 wl_113 vdd gnd cell_6t
Xbit_r114_c5 bl_5 br_5 wl_114 vdd gnd cell_6t
Xbit_r115_c5 bl_5 br_5 wl_115 vdd gnd cell_6t
Xbit_r116_c5 bl_5 br_5 wl_116 vdd gnd cell_6t
Xbit_r117_c5 bl_5 br_5 wl_117 vdd gnd cell_6t
Xbit_r118_c5 bl_5 br_5 wl_118 vdd gnd cell_6t
Xbit_r119_c5 bl_5 br_5 wl_119 vdd gnd cell_6t
Xbit_r120_c5 bl_5 br_5 wl_120 vdd gnd cell_6t
Xbit_r121_c5 bl_5 br_5 wl_121 vdd gnd cell_6t
Xbit_r122_c5 bl_5 br_5 wl_122 vdd gnd cell_6t
Xbit_r123_c5 bl_5 br_5 wl_123 vdd gnd cell_6t
Xbit_r124_c5 bl_5 br_5 wl_124 vdd gnd cell_6t
Xbit_r125_c5 bl_5 br_5 wl_125 vdd gnd cell_6t
Xbit_r126_c5 bl_5 br_5 wl_126 vdd gnd cell_6t
Xbit_r127_c5 bl_5 br_5 wl_127 vdd gnd cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd cell_6t
Xbit_r1_c6 bl_6 br_6 wl_1 vdd gnd cell_6t
Xbit_r2_c6 bl_6 br_6 wl_2 vdd gnd cell_6t
Xbit_r3_c6 bl_6 br_6 wl_3 vdd gnd cell_6t
Xbit_r4_c6 bl_6 br_6 wl_4 vdd gnd cell_6t
Xbit_r5_c6 bl_6 br_6 wl_5 vdd gnd cell_6t
Xbit_r6_c6 bl_6 br_6 wl_6 vdd gnd cell_6t
Xbit_r7_c6 bl_6 br_6 wl_7 vdd gnd cell_6t
Xbit_r8_c6 bl_6 br_6 wl_8 vdd gnd cell_6t
Xbit_r9_c6 bl_6 br_6 wl_9 vdd gnd cell_6t
Xbit_r10_c6 bl_6 br_6 wl_10 vdd gnd cell_6t
Xbit_r11_c6 bl_6 br_6 wl_11 vdd gnd cell_6t
Xbit_r12_c6 bl_6 br_6 wl_12 vdd gnd cell_6t
Xbit_r13_c6 bl_6 br_6 wl_13 vdd gnd cell_6t
Xbit_r14_c6 bl_6 br_6 wl_14 vdd gnd cell_6t
Xbit_r15_c6 bl_6 br_6 wl_15 vdd gnd cell_6t
Xbit_r16_c6 bl_6 br_6 wl_16 vdd gnd cell_6t
Xbit_r17_c6 bl_6 br_6 wl_17 vdd gnd cell_6t
Xbit_r18_c6 bl_6 br_6 wl_18 vdd gnd cell_6t
Xbit_r19_c6 bl_6 br_6 wl_19 vdd gnd cell_6t
Xbit_r20_c6 bl_6 br_6 wl_20 vdd gnd cell_6t
Xbit_r21_c6 bl_6 br_6 wl_21 vdd gnd cell_6t
Xbit_r22_c6 bl_6 br_6 wl_22 vdd gnd cell_6t
Xbit_r23_c6 bl_6 br_6 wl_23 vdd gnd cell_6t
Xbit_r24_c6 bl_6 br_6 wl_24 vdd gnd cell_6t
Xbit_r25_c6 bl_6 br_6 wl_25 vdd gnd cell_6t
Xbit_r26_c6 bl_6 br_6 wl_26 vdd gnd cell_6t
Xbit_r27_c6 bl_6 br_6 wl_27 vdd gnd cell_6t
Xbit_r28_c6 bl_6 br_6 wl_28 vdd gnd cell_6t
Xbit_r29_c6 bl_6 br_6 wl_29 vdd gnd cell_6t
Xbit_r30_c6 bl_6 br_6 wl_30 vdd gnd cell_6t
Xbit_r31_c6 bl_6 br_6 wl_31 vdd gnd cell_6t
Xbit_r32_c6 bl_6 br_6 wl_32 vdd gnd cell_6t
Xbit_r33_c6 bl_6 br_6 wl_33 vdd gnd cell_6t
Xbit_r34_c6 bl_6 br_6 wl_34 vdd gnd cell_6t
Xbit_r35_c6 bl_6 br_6 wl_35 vdd gnd cell_6t
Xbit_r36_c6 bl_6 br_6 wl_36 vdd gnd cell_6t
Xbit_r37_c6 bl_6 br_6 wl_37 vdd gnd cell_6t
Xbit_r38_c6 bl_6 br_6 wl_38 vdd gnd cell_6t
Xbit_r39_c6 bl_6 br_6 wl_39 vdd gnd cell_6t
Xbit_r40_c6 bl_6 br_6 wl_40 vdd gnd cell_6t
Xbit_r41_c6 bl_6 br_6 wl_41 vdd gnd cell_6t
Xbit_r42_c6 bl_6 br_6 wl_42 vdd gnd cell_6t
Xbit_r43_c6 bl_6 br_6 wl_43 vdd gnd cell_6t
Xbit_r44_c6 bl_6 br_6 wl_44 vdd gnd cell_6t
Xbit_r45_c6 bl_6 br_6 wl_45 vdd gnd cell_6t
Xbit_r46_c6 bl_6 br_6 wl_46 vdd gnd cell_6t
Xbit_r47_c6 bl_6 br_6 wl_47 vdd gnd cell_6t
Xbit_r48_c6 bl_6 br_6 wl_48 vdd gnd cell_6t
Xbit_r49_c6 bl_6 br_6 wl_49 vdd gnd cell_6t
Xbit_r50_c6 bl_6 br_6 wl_50 vdd gnd cell_6t
Xbit_r51_c6 bl_6 br_6 wl_51 vdd gnd cell_6t
Xbit_r52_c6 bl_6 br_6 wl_52 vdd gnd cell_6t
Xbit_r53_c6 bl_6 br_6 wl_53 vdd gnd cell_6t
Xbit_r54_c6 bl_6 br_6 wl_54 vdd gnd cell_6t
Xbit_r55_c6 bl_6 br_6 wl_55 vdd gnd cell_6t
Xbit_r56_c6 bl_6 br_6 wl_56 vdd gnd cell_6t
Xbit_r57_c6 bl_6 br_6 wl_57 vdd gnd cell_6t
Xbit_r58_c6 bl_6 br_6 wl_58 vdd gnd cell_6t
Xbit_r59_c6 bl_6 br_6 wl_59 vdd gnd cell_6t
Xbit_r60_c6 bl_6 br_6 wl_60 vdd gnd cell_6t
Xbit_r61_c6 bl_6 br_6 wl_61 vdd gnd cell_6t
Xbit_r62_c6 bl_6 br_6 wl_62 vdd gnd cell_6t
Xbit_r63_c6 bl_6 br_6 wl_63 vdd gnd cell_6t
Xbit_r64_c6 bl_6 br_6 wl_64 vdd gnd cell_6t
Xbit_r65_c6 bl_6 br_6 wl_65 vdd gnd cell_6t
Xbit_r66_c6 bl_6 br_6 wl_66 vdd gnd cell_6t
Xbit_r67_c6 bl_6 br_6 wl_67 vdd gnd cell_6t
Xbit_r68_c6 bl_6 br_6 wl_68 vdd gnd cell_6t
Xbit_r69_c6 bl_6 br_6 wl_69 vdd gnd cell_6t
Xbit_r70_c6 bl_6 br_6 wl_70 vdd gnd cell_6t
Xbit_r71_c6 bl_6 br_6 wl_71 vdd gnd cell_6t
Xbit_r72_c6 bl_6 br_6 wl_72 vdd gnd cell_6t
Xbit_r73_c6 bl_6 br_6 wl_73 vdd gnd cell_6t
Xbit_r74_c6 bl_6 br_6 wl_74 vdd gnd cell_6t
Xbit_r75_c6 bl_6 br_6 wl_75 vdd gnd cell_6t
Xbit_r76_c6 bl_6 br_6 wl_76 vdd gnd cell_6t
Xbit_r77_c6 bl_6 br_6 wl_77 vdd gnd cell_6t
Xbit_r78_c6 bl_6 br_6 wl_78 vdd gnd cell_6t
Xbit_r79_c6 bl_6 br_6 wl_79 vdd gnd cell_6t
Xbit_r80_c6 bl_6 br_6 wl_80 vdd gnd cell_6t
Xbit_r81_c6 bl_6 br_6 wl_81 vdd gnd cell_6t
Xbit_r82_c6 bl_6 br_6 wl_82 vdd gnd cell_6t
Xbit_r83_c6 bl_6 br_6 wl_83 vdd gnd cell_6t
Xbit_r84_c6 bl_6 br_6 wl_84 vdd gnd cell_6t
Xbit_r85_c6 bl_6 br_6 wl_85 vdd gnd cell_6t
Xbit_r86_c6 bl_6 br_6 wl_86 vdd gnd cell_6t
Xbit_r87_c6 bl_6 br_6 wl_87 vdd gnd cell_6t
Xbit_r88_c6 bl_6 br_6 wl_88 vdd gnd cell_6t
Xbit_r89_c6 bl_6 br_6 wl_89 vdd gnd cell_6t
Xbit_r90_c6 bl_6 br_6 wl_90 vdd gnd cell_6t
Xbit_r91_c6 bl_6 br_6 wl_91 vdd gnd cell_6t
Xbit_r92_c6 bl_6 br_6 wl_92 vdd gnd cell_6t
Xbit_r93_c6 bl_6 br_6 wl_93 vdd gnd cell_6t
Xbit_r94_c6 bl_6 br_6 wl_94 vdd gnd cell_6t
Xbit_r95_c6 bl_6 br_6 wl_95 vdd gnd cell_6t
Xbit_r96_c6 bl_6 br_6 wl_96 vdd gnd cell_6t
Xbit_r97_c6 bl_6 br_6 wl_97 vdd gnd cell_6t
Xbit_r98_c6 bl_6 br_6 wl_98 vdd gnd cell_6t
Xbit_r99_c6 bl_6 br_6 wl_99 vdd gnd cell_6t
Xbit_r100_c6 bl_6 br_6 wl_100 vdd gnd cell_6t
Xbit_r101_c6 bl_6 br_6 wl_101 vdd gnd cell_6t
Xbit_r102_c6 bl_6 br_6 wl_102 vdd gnd cell_6t
Xbit_r103_c6 bl_6 br_6 wl_103 vdd gnd cell_6t
Xbit_r104_c6 bl_6 br_6 wl_104 vdd gnd cell_6t
Xbit_r105_c6 bl_6 br_6 wl_105 vdd gnd cell_6t
Xbit_r106_c6 bl_6 br_6 wl_106 vdd gnd cell_6t
Xbit_r107_c6 bl_6 br_6 wl_107 vdd gnd cell_6t
Xbit_r108_c6 bl_6 br_6 wl_108 vdd gnd cell_6t
Xbit_r109_c6 bl_6 br_6 wl_109 vdd gnd cell_6t
Xbit_r110_c6 bl_6 br_6 wl_110 vdd gnd cell_6t
Xbit_r111_c6 bl_6 br_6 wl_111 vdd gnd cell_6t
Xbit_r112_c6 bl_6 br_6 wl_112 vdd gnd cell_6t
Xbit_r113_c6 bl_6 br_6 wl_113 vdd gnd cell_6t
Xbit_r114_c6 bl_6 br_6 wl_114 vdd gnd cell_6t
Xbit_r115_c6 bl_6 br_6 wl_115 vdd gnd cell_6t
Xbit_r116_c6 bl_6 br_6 wl_116 vdd gnd cell_6t
Xbit_r117_c6 bl_6 br_6 wl_117 vdd gnd cell_6t
Xbit_r118_c6 bl_6 br_6 wl_118 vdd gnd cell_6t
Xbit_r119_c6 bl_6 br_6 wl_119 vdd gnd cell_6t
Xbit_r120_c6 bl_6 br_6 wl_120 vdd gnd cell_6t
Xbit_r121_c6 bl_6 br_6 wl_121 vdd gnd cell_6t
Xbit_r122_c6 bl_6 br_6 wl_122 vdd gnd cell_6t
Xbit_r123_c6 bl_6 br_6 wl_123 vdd gnd cell_6t
Xbit_r124_c6 bl_6 br_6 wl_124 vdd gnd cell_6t
Xbit_r125_c6 bl_6 br_6 wl_125 vdd gnd cell_6t
Xbit_r126_c6 bl_6 br_6 wl_126 vdd gnd cell_6t
Xbit_r127_c6 bl_6 br_6 wl_127 vdd gnd cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd cell_6t
Xbit_r1_c7 bl_7 br_7 wl_1 vdd gnd cell_6t
Xbit_r2_c7 bl_7 br_7 wl_2 vdd gnd cell_6t
Xbit_r3_c7 bl_7 br_7 wl_3 vdd gnd cell_6t
Xbit_r4_c7 bl_7 br_7 wl_4 vdd gnd cell_6t
Xbit_r5_c7 bl_7 br_7 wl_5 vdd gnd cell_6t
Xbit_r6_c7 bl_7 br_7 wl_6 vdd gnd cell_6t
Xbit_r7_c7 bl_7 br_7 wl_7 vdd gnd cell_6t
Xbit_r8_c7 bl_7 br_7 wl_8 vdd gnd cell_6t
Xbit_r9_c7 bl_7 br_7 wl_9 vdd gnd cell_6t
Xbit_r10_c7 bl_7 br_7 wl_10 vdd gnd cell_6t
Xbit_r11_c7 bl_7 br_7 wl_11 vdd gnd cell_6t
Xbit_r12_c7 bl_7 br_7 wl_12 vdd gnd cell_6t
Xbit_r13_c7 bl_7 br_7 wl_13 vdd gnd cell_6t
Xbit_r14_c7 bl_7 br_7 wl_14 vdd gnd cell_6t
Xbit_r15_c7 bl_7 br_7 wl_15 vdd gnd cell_6t
Xbit_r16_c7 bl_7 br_7 wl_16 vdd gnd cell_6t
Xbit_r17_c7 bl_7 br_7 wl_17 vdd gnd cell_6t
Xbit_r18_c7 bl_7 br_7 wl_18 vdd gnd cell_6t
Xbit_r19_c7 bl_7 br_7 wl_19 vdd gnd cell_6t
Xbit_r20_c7 bl_7 br_7 wl_20 vdd gnd cell_6t
Xbit_r21_c7 bl_7 br_7 wl_21 vdd gnd cell_6t
Xbit_r22_c7 bl_7 br_7 wl_22 vdd gnd cell_6t
Xbit_r23_c7 bl_7 br_7 wl_23 vdd gnd cell_6t
Xbit_r24_c7 bl_7 br_7 wl_24 vdd gnd cell_6t
Xbit_r25_c7 bl_7 br_7 wl_25 vdd gnd cell_6t
Xbit_r26_c7 bl_7 br_7 wl_26 vdd gnd cell_6t
Xbit_r27_c7 bl_7 br_7 wl_27 vdd gnd cell_6t
Xbit_r28_c7 bl_7 br_7 wl_28 vdd gnd cell_6t
Xbit_r29_c7 bl_7 br_7 wl_29 vdd gnd cell_6t
Xbit_r30_c7 bl_7 br_7 wl_30 vdd gnd cell_6t
Xbit_r31_c7 bl_7 br_7 wl_31 vdd gnd cell_6t
Xbit_r32_c7 bl_7 br_7 wl_32 vdd gnd cell_6t
Xbit_r33_c7 bl_7 br_7 wl_33 vdd gnd cell_6t
Xbit_r34_c7 bl_7 br_7 wl_34 vdd gnd cell_6t
Xbit_r35_c7 bl_7 br_7 wl_35 vdd gnd cell_6t
Xbit_r36_c7 bl_7 br_7 wl_36 vdd gnd cell_6t
Xbit_r37_c7 bl_7 br_7 wl_37 vdd gnd cell_6t
Xbit_r38_c7 bl_7 br_7 wl_38 vdd gnd cell_6t
Xbit_r39_c7 bl_7 br_7 wl_39 vdd gnd cell_6t
Xbit_r40_c7 bl_7 br_7 wl_40 vdd gnd cell_6t
Xbit_r41_c7 bl_7 br_7 wl_41 vdd gnd cell_6t
Xbit_r42_c7 bl_7 br_7 wl_42 vdd gnd cell_6t
Xbit_r43_c7 bl_7 br_7 wl_43 vdd gnd cell_6t
Xbit_r44_c7 bl_7 br_7 wl_44 vdd gnd cell_6t
Xbit_r45_c7 bl_7 br_7 wl_45 vdd gnd cell_6t
Xbit_r46_c7 bl_7 br_7 wl_46 vdd gnd cell_6t
Xbit_r47_c7 bl_7 br_7 wl_47 vdd gnd cell_6t
Xbit_r48_c7 bl_7 br_7 wl_48 vdd gnd cell_6t
Xbit_r49_c7 bl_7 br_7 wl_49 vdd gnd cell_6t
Xbit_r50_c7 bl_7 br_7 wl_50 vdd gnd cell_6t
Xbit_r51_c7 bl_7 br_7 wl_51 vdd gnd cell_6t
Xbit_r52_c7 bl_7 br_7 wl_52 vdd gnd cell_6t
Xbit_r53_c7 bl_7 br_7 wl_53 vdd gnd cell_6t
Xbit_r54_c7 bl_7 br_7 wl_54 vdd gnd cell_6t
Xbit_r55_c7 bl_7 br_7 wl_55 vdd gnd cell_6t
Xbit_r56_c7 bl_7 br_7 wl_56 vdd gnd cell_6t
Xbit_r57_c7 bl_7 br_7 wl_57 vdd gnd cell_6t
Xbit_r58_c7 bl_7 br_7 wl_58 vdd gnd cell_6t
Xbit_r59_c7 bl_7 br_7 wl_59 vdd gnd cell_6t
Xbit_r60_c7 bl_7 br_7 wl_60 vdd gnd cell_6t
Xbit_r61_c7 bl_7 br_7 wl_61 vdd gnd cell_6t
Xbit_r62_c7 bl_7 br_7 wl_62 vdd gnd cell_6t
Xbit_r63_c7 bl_7 br_7 wl_63 vdd gnd cell_6t
Xbit_r64_c7 bl_7 br_7 wl_64 vdd gnd cell_6t
Xbit_r65_c7 bl_7 br_7 wl_65 vdd gnd cell_6t
Xbit_r66_c7 bl_7 br_7 wl_66 vdd gnd cell_6t
Xbit_r67_c7 bl_7 br_7 wl_67 vdd gnd cell_6t
Xbit_r68_c7 bl_7 br_7 wl_68 vdd gnd cell_6t
Xbit_r69_c7 bl_7 br_7 wl_69 vdd gnd cell_6t
Xbit_r70_c7 bl_7 br_7 wl_70 vdd gnd cell_6t
Xbit_r71_c7 bl_7 br_7 wl_71 vdd gnd cell_6t
Xbit_r72_c7 bl_7 br_7 wl_72 vdd gnd cell_6t
Xbit_r73_c7 bl_7 br_7 wl_73 vdd gnd cell_6t
Xbit_r74_c7 bl_7 br_7 wl_74 vdd gnd cell_6t
Xbit_r75_c7 bl_7 br_7 wl_75 vdd gnd cell_6t
Xbit_r76_c7 bl_7 br_7 wl_76 vdd gnd cell_6t
Xbit_r77_c7 bl_7 br_7 wl_77 vdd gnd cell_6t
Xbit_r78_c7 bl_7 br_7 wl_78 vdd gnd cell_6t
Xbit_r79_c7 bl_7 br_7 wl_79 vdd gnd cell_6t
Xbit_r80_c7 bl_7 br_7 wl_80 vdd gnd cell_6t
Xbit_r81_c7 bl_7 br_7 wl_81 vdd gnd cell_6t
Xbit_r82_c7 bl_7 br_7 wl_82 vdd gnd cell_6t
Xbit_r83_c7 bl_7 br_7 wl_83 vdd gnd cell_6t
Xbit_r84_c7 bl_7 br_7 wl_84 vdd gnd cell_6t
Xbit_r85_c7 bl_7 br_7 wl_85 vdd gnd cell_6t
Xbit_r86_c7 bl_7 br_7 wl_86 vdd gnd cell_6t
Xbit_r87_c7 bl_7 br_7 wl_87 vdd gnd cell_6t
Xbit_r88_c7 bl_7 br_7 wl_88 vdd gnd cell_6t
Xbit_r89_c7 bl_7 br_7 wl_89 vdd gnd cell_6t
Xbit_r90_c7 bl_7 br_7 wl_90 vdd gnd cell_6t
Xbit_r91_c7 bl_7 br_7 wl_91 vdd gnd cell_6t
Xbit_r92_c7 bl_7 br_7 wl_92 vdd gnd cell_6t
Xbit_r93_c7 bl_7 br_7 wl_93 vdd gnd cell_6t
Xbit_r94_c7 bl_7 br_7 wl_94 vdd gnd cell_6t
Xbit_r95_c7 bl_7 br_7 wl_95 vdd gnd cell_6t
Xbit_r96_c7 bl_7 br_7 wl_96 vdd gnd cell_6t
Xbit_r97_c7 bl_7 br_7 wl_97 vdd gnd cell_6t
Xbit_r98_c7 bl_7 br_7 wl_98 vdd gnd cell_6t
Xbit_r99_c7 bl_7 br_7 wl_99 vdd gnd cell_6t
Xbit_r100_c7 bl_7 br_7 wl_100 vdd gnd cell_6t
Xbit_r101_c7 bl_7 br_7 wl_101 vdd gnd cell_6t
Xbit_r102_c7 bl_7 br_7 wl_102 vdd gnd cell_6t
Xbit_r103_c7 bl_7 br_7 wl_103 vdd gnd cell_6t
Xbit_r104_c7 bl_7 br_7 wl_104 vdd gnd cell_6t
Xbit_r105_c7 bl_7 br_7 wl_105 vdd gnd cell_6t
Xbit_r106_c7 bl_7 br_7 wl_106 vdd gnd cell_6t
Xbit_r107_c7 bl_7 br_7 wl_107 vdd gnd cell_6t
Xbit_r108_c7 bl_7 br_7 wl_108 vdd gnd cell_6t
Xbit_r109_c7 bl_7 br_7 wl_109 vdd gnd cell_6t
Xbit_r110_c7 bl_7 br_7 wl_110 vdd gnd cell_6t
Xbit_r111_c7 bl_7 br_7 wl_111 vdd gnd cell_6t
Xbit_r112_c7 bl_7 br_7 wl_112 vdd gnd cell_6t
Xbit_r113_c7 bl_7 br_7 wl_113 vdd gnd cell_6t
Xbit_r114_c7 bl_7 br_7 wl_114 vdd gnd cell_6t
Xbit_r115_c7 bl_7 br_7 wl_115 vdd gnd cell_6t
Xbit_r116_c7 bl_7 br_7 wl_116 vdd gnd cell_6t
Xbit_r117_c7 bl_7 br_7 wl_117 vdd gnd cell_6t
Xbit_r118_c7 bl_7 br_7 wl_118 vdd gnd cell_6t
Xbit_r119_c7 bl_7 br_7 wl_119 vdd gnd cell_6t
Xbit_r120_c7 bl_7 br_7 wl_120 vdd gnd cell_6t
Xbit_r121_c7 bl_7 br_7 wl_121 vdd gnd cell_6t
Xbit_r122_c7 bl_7 br_7 wl_122 vdd gnd cell_6t
Xbit_r123_c7 bl_7 br_7 wl_123 vdd gnd cell_6t
Xbit_r124_c7 bl_7 br_7 wl_124 vdd gnd cell_6t
Xbit_r125_c7 bl_7 br_7 wl_125 vdd gnd cell_6t
Xbit_r126_c7 bl_7 br_7 wl_126 vdd gnd cell_6t
Xbit_r127_c7 bl_7 br_7 wl_127 vdd gnd cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd cell_6t
Xbit_r1_c8 bl_8 br_8 wl_1 vdd gnd cell_6t
Xbit_r2_c8 bl_8 br_8 wl_2 vdd gnd cell_6t
Xbit_r3_c8 bl_8 br_8 wl_3 vdd gnd cell_6t
Xbit_r4_c8 bl_8 br_8 wl_4 vdd gnd cell_6t
Xbit_r5_c8 bl_8 br_8 wl_5 vdd gnd cell_6t
Xbit_r6_c8 bl_8 br_8 wl_6 vdd gnd cell_6t
Xbit_r7_c8 bl_8 br_8 wl_7 vdd gnd cell_6t
Xbit_r8_c8 bl_8 br_8 wl_8 vdd gnd cell_6t
Xbit_r9_c8 bl_8 br_8 wl_9 vdd gnd cell_6t
Xbit_r10_c8 bl_8 br_8 wl_10 vdd gnd cell_6t
Xbit_r11_c8 bl_8 br_8 wl_11 vdd gnd cell_6t
Xbit_r12_c8 bl_8 br_8 wl_12 vdd gnd cell_6t
Xbit_r13_c8 bl_8 br_8 wl_13 vdd gnd cell_6t
Xbit_r14_c8 bl_8 br_8 wl_14 vdd gnd cell_6t
Xbit_r15_c8 bl_8 br_8 wl_15 vdd gnd cell_6t
Xbit_r16_c8 bl_8 br_8 wl_16 vdd gnd cell_6t
Xbit_r17_c8 bl_8 br_8 wl_17 vdd gnd cell_6t
Xbit_r18_c8 bl_8 br_8 wl_18 vdd gnd cell_6t
Xbit_r19_c8 bl_8 br_8 wl_19 vdd gnd cell_6t
Xbit_r20_c8 bl_8 br_8 wl_20 vdd gnd cell_6t
Xbit_r21_c8 bl_8 br_8 wl_21 vdd gnd cell_6t
Xbit_r22_c8 bl_8 br_8 wl_22 vdd gnd cell_6t
Xbit_r23_c8 bl_8 br_8 wl_23 vdd gnd cell_6t
Xbit_r24_c8 bl_8 br_8 wl_24 vdd gnd cell_6t
Xbit_r25_c8 bl_8 br_8 wl_25 vdd gnd cell_6t
Xbit_r26_c8 bl_8 br_8 wl_26 vdd gnd cell_6t
Xbit_r27_c8 bl_8 br_8 wl_27 vdd gnd cell_6t
Xbit_r28_c8 bl_8 br_8 wl_28 vdd gnd cell_6t
Xbit_r29_c8 bl_8 br_8 wl_29 vdd gnd cell_6t
Xbit_r30_c8 bl_8 br_8 wl_30 vdd gnd cell_6t
Xbit_r31_c8 bl_8 br_8 wl_31 vdd gnd cell_6t
Xbit_r32_c8 bl_8 br_8 wl_32 vdd gnd cell_6t
Xbit_r33_c8 bl_8 br_8 wl_33 vdd gnd cell_6t
Xbit_r34_c8 bl_8 br_8 wl_34 vdd gnd cell_6t
Xbit_r35_c8 bl_8 br_8 wl_35 vdd gnd cell_6t
Xbit_r36_c8 bl_8 br_8 wl_36 vdd gnd cell_6t
Xbit_r37_c8 bl_8 br_8 wl_37 vdd gnd cell_6t
Xbit_r38_c8 bl_8 br_8 wl_38 vdd gnd cell_6t
Xbit_r39_c8 bl_8 br_8 wl_39 vdd gnd cell_6t
Xbit_r40_c8 bl_8 br_8 wl_40 vdd gnd cell_6t
Xbit_r41_c8 bl_8 br_8 wl_41 vdd gnd cell_6t
Xbit_r42_c8 bl_8 br_8 wl_42 vdd gnd cell_6t
Xbit_r43_c8 bl_8 br_8 wl_43 vdd gnd cell_6t
Xbit_r44_c8 bl_8 br_8 wl_44 vdd gnd cell_6t
Xbit_r45_c8 bl_8 br_8 wl_45 vdd gnd cell_6t
Xbit_r46_c8 bl_8 br_8 wl_46 vdd gnd cell_6t
Xbit_r47_c8 bl_8 br_8 wl_47 vdd gnd cell_6t
Xbit_r48_c8 bl_8 br_8 wl_48 vdd gnd cell_6t
Xbit_r49_c8 bl_8 br_8 wl_49 vdd gnd cell_6t
Xbit_r50_c8 bl_8 br_8 wl_50 vdd gnd cell_6t
Xbit_r51_c8 bl_8 br_8 wl_51 vdd gnd cell_6t
Xbit_r52_c8 bl_8 br_8 wl_52 vdd gnd cell_6t
Xbit_r53_c8 bl_8 br_8 wl_53 vdd gnd cell_6t
Xbit_r54_c8 bl_8 br_8 wl_54 vdd gnd cell_6t
Xbit_r55_c8 bl_8 br_8 wl_55 vdd gnd cell_6t
Xbit_r56_c8 bl_8 br_8 wl_56 vdd gnd cell_6t
Xbit_r57_c8 bl_8 br_8 wl_57 vdd gnd cell_6t
Xbit_r58_c8 bl_8 br_8 wl_58 vdd gnd cell_6t
Xbit_r59_c8 bl_8 br_8 wl_59 vdd gnd cell_6t
Xbit_r60_c8 bl_8 br_8 wl_60 vdd gnd cell_6t
Xbit_r61_c8 bl_8 br_8 wl_61 vdd gnd cell_6t
Xbit_r62_c8 bl_8 br_8 wl_62 vdd gnd cell_6t
Xbit_r63_c8 bl_8 br_8 wl_63 vdd gnd cell_6t
Xbit_r64_c8 bl_8 br_8 wl_64 vdd gnd cell_6t
Xbit_r65_c8 bl_8 br_8 wl_65 vdd gnd cell_6t
Xbit_r66_c8 bl_8 br_8 wl_66 vdd gnd cell_6t
Xbit_r67_c8 bl_8 br_8 wl_67 vdd gnd cell_6t
Xbit_r68_c8 bl_8 br_8 wl_68 vdd gnd cell_6t
Xbit_r69_c8 bl_8 br_8 wl_69 vdd gnd cell_6t
Xbit_r70_c8 bl_8 br_8 wl_70 vdd gnd cell_6t
Xbit_r71_c8 bl_8 br_8 wl_71 vdd gnd cell_6t
Xbit_r72_c8 bl_8 br_8 wl_72 vdd gnd cell_6t
Xbit_r73_c8 bl_8 br_8 wl_73 vdd gnd cell_6t
Xbit_r74_c8 bl_8 br_8 wl_74 vdd gnd cell_6t
Xbit_r75_c8 bl_8 br_8 wl_75 vdd gnd cell_6t
Xbit_r76_c8 bl_8 br_8 wl_76 vdd gnd cell_6t
Xbit_r77_c8 bl_8 br_8 wl_77 vdd gnd cell_6t
Xbit_r78_c8 bl_8 br_8 wl_78 vdd gnd cell_6t
Xbit_r79_c8 bl_8 br_8 wl_79 vdd gnd cell_6t
Xbit_r80_c8 bl_8 br_8 wl_80 vdd gnd cell_6t
Xbit_r81_c8 bl_8 br_8 wl_81 vdd gnd cell_6t
Xbit_r82_c8 bl_8 br_8 wl_82 vdd gnd cell_6t
Xbit_r83_c8 bl_8 br_8 wl_83 vdd gnd cell_6t
Xbit_r84_c8 bl_8 br_8 wl_84 vdd gnd cell_6t
Xbit_r85_c8 bl_8 br_8 wl_85 vdd gnd cell_6t
Xbit_r86_c8 bl_8 br_8 wl_86 vdd gnd cell_6t
Xbit_r87_c8 bl_8 br_8 wl_87 vdd gnd cell_6t
Xbit_r88_c8 bl_8 br_8 wl_88 vdd gnd cell_6t
Xbit_r89_c8 bl_8 br_8 wl_89 vdd gnd cell_6t
Xbit_r90_c8 bl_8 br_8 wl_90 vdd gnd cell_6t
Xbit_r91_c8 bl_8 br_8 wl_91 vdd gnd cell_6t
Xbit_r92_c8 bl_8 br_8 wl_92 vdd gnd cell_6t
Xbit_r93_c8 bl_8 br_8 wl_93 vdd gnd cell_6t
Xbit_r94_c8 bl_8 br_8 wl_94 vdd gnd cell_6t
Xbit_r95_c8 bl_8 br_8 wl_95 vdd gnd cell_6t
Xbit_r96_c8 bl_8 br_8 wl_96 vdd gnd cell_6t
Xbit_r97_c8 bl_8 br_8 wl_97 vdd gnd cell_6t
Xbit_r98_c8 bl_8 br_8 wl_98 vdd gnd cell_6t
Xbit_r99_c8 bl_8 br_8 wl_99 vdd gnd cell_6t
Xbit_r100_c8 bl_8 br_8 wl_100 vdd gnd cell_6t
Xbit_r101_c8 bl_8 br_8 wl_101 vdd gnd cell_6t
Xbit_r102_c8 bl_8 br_8 wl_102 vdd gnd cell_6t
Xbit_r103_c8 bl_8 br_8 wl_103 vdd gnd cell_6t
Xbit_r104_c8 bl_8 br_8 wl_104 vdd gnd cell_6t
Xbit_r105_c8 bl_8 br_8 wl_105 vdd gnd cell_6t
Xbit_r106_c8 bl_8 br_8 wl_106 vdd gnd cell_6t
Xbit_r107_c8 bl_8 br_8 wl_107 vdd gnd cell_6t
Xbit_r108_c8 bl_8 br_8 wl_108 vdd gnd cell_6t
Xbit_r109_c8 bl_8 br_8 wl_109 vdd gnd cell_6t
Xbit_r110_c8 bl_8 br_8 wl_110 vdd gnd cell_6t
Xbit_r111_c8 bl_8 br_8 wl_111 vdd gnd cell_6t
Xbit_r112_c8 bl_8 br_8 wl_112 vdd gnd cell_6t
Xbit_r113_c8 bl_8 br_8 wl_113 vdd gnd cell_6t
Xbit_r114_c8 bl_8 br_8 wl_114 vdd gnd cell_6t
Xbit_r115_c8 bl_8 br_8 wl_115 vdd gnd cell_6t
Xbit_r116_c8 bl_8 br_8 wl_116 vdd gnd cell_6t
Xbit_r117_c8 bl_8 br_8 wl_117 vdd gnd cell_6t
Xbit_r118_c8 bl_8 br_8 wl_118 vdd gnd cell_6t
Xbit_r119_c8 bl_8 br_8 wl_119 vdd gnd cell_6t
Xbit_r120_c8 bl_8 br_8 wl_120 vdd gnd cell_6t
Xbit_r121_c8 bl_8 br_8 wl_121 vdd gnd cell_6t
Xbit_r122_c8 bl_8 br_8 wl_122 vdd gnd cell_6t
Xbit_r123_c8 bl_8 br_8 wl_123 vdd gnd cell_6t
Xbit_r124_c8 bl_8 br_8 wl_124 vdd gnd cell_6t
Xbit_r125_c8 bl_8 br_8 wl_125 vdd gnd cell_6t
Xbit_r126_c8 bl_8 br_8 wl_126 vdd gnd cell_6t
Xbit_r127_c8 bl_8 br_8 wl_127 vdd gnd cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd cell_6t
Xbit_r1_c9 bl_9 br_9 wl_1 vdd gnd cell_6t
Xbit_r2_c9 bl_9 br_9 wl_2 vdd gnd cell_6t
Xbit_r3_c9 bl_9 br_9 wl_3 vdd gnd cell_6t
Xbit_r4_c9 bl_9 br_9 wl_4 vdd gnd cell_6t
Xbit_r5_c9 bl_9 br_9 wl_5 vdd gnd cell_6t
Xbit_r6_c9 bl_9 br_9 wl_6 vdd gnd cell_6t
Xbit_r7_c9 bl_9 br_9 wl_7 vdd gnd cell_6t
Xbit_r8_c9 bl_9 br_9 wl_8 vdd gnd cell_6t
Xbit_r9_c9 bl_9 br_9 wl_9 vdd gnd cell_6t
Xbit_r10_c9 bl_9 br_9 wl_10 vdd gnd cell_6t
Xbit_r11_c9 bl_9 br_9 wl_11 vdd gnd cell_6t
Xbit_r12_c9 bl_9 br_9 wl_12 vdd gnd cell_6t
Xbit_r13_c9 bl_9 br_9 wl_13 vdd gnd cell_6t
Xbit_r14_c9 bl_9 br_9 wl_14 vdd gnd cell_6t
Xbit_r15_c9 bl_9 br_9 wl_15 vdd gnd cell_6t
Xbit_r16_c9 bl_9 br_9 wl_16 vdd gnd cell_6t
Xbit_r17_c9 bl_9 br_9 wl_17 vdd gnd cell_6t
Xbit_r18_c9 bl_9 br_9 wl_18 vdd gnd cell_6t
Xbit_r19_c9 bl_9 br_9 wl_19 vdd gnd cell_6t
Xbit_r20_c9 bl_9 br_9 wl_20 vdd gnd cell_6t
Xbit_r21_c9 bl_9 br_9 wl_21 vdd gnd cell_6t
Xbit_r22_c9 bl_9 br_9 wl_22 vdd gnd cell_6t
Xbit_r23_c9 bl_9 br_9 wl_23 vdd gnd cell_6t
Xbit_r24_c9 bl_9 br_9 wl_24 vdd gnd cell_6t
Xbit_r25_c9 bl_9 br_9 wl_25 vdd gnd cell_6t
Xbit_r26_c9 bl_9 br_9 wl_26 vdd gnd cell_6t
Xbit_r27_c9 bl_9 br_9 wl_27 vdd gnd cell_6t
Xbit_r28_c9 bl_9 br_9 wl_28 vdd gnd cell_6t
Xbit_r29_c9 bl_9 br_9 wl_29 vdd gnd cell_6t
Xbit_r30_c9 bl_9 br_9 wl_30 vdd gnd cell_6t
Xbit_r31_c9 bl_9 br_9 wl_31 vdd gnd cell_6t
Xbit_r32_c9 bl_9 br_9 wl_32 vdd gnd cell_6t
Xbit_r33_c9 bl_9 br_9 wl_33 vdd gnd cell_6t
Xbit_r34_c9 bl_9 br_9 wl_34 vdd gnd cell_6t
Xbit_r35_c9 bl_9 br_9 wl_35 vdd gnd cell_6t
Xbit_r36_c9 bl_9 br_9 wl_36 vdd gnd cell_6t
Xbit_r37_c9 bl_9 br_9 wl_37 vdd gnd cell_6t
Xbit_r38_c9 bl_9 br_9 wl_38 vdd gnd cell_6t
Xbit_r39_c9 bl_9 br_9 wl_39 vdd gnd cell_6t
Xbit_r40_c9 bl_9 br_9 wl_40 vdd gnd cell_6t
Xbit_r41_c9 bl_9 br_9 wl_41 vdd gnd cell_6t
Xbit_r42_c9 bl_9 br_9 wl_42 vdd gnd cell_6t
Xbit_r43_c9 bl_9 br_9 wl_43 vdd gnd cell_6t
Xbit_r44_c9 bl_9 br_9 wl_44 vdd gnd cell_6t
Xbit_r45_c9 bl_9 br_9 wl_45 vdd gnd cell_6t
Xbit_r46_c9 bl_9 br_9 wl_46 vdd gnd cell_6t
Xbit_r47_c9 bl_9 br_9 wl_47 vdd gnd cell_6t
Xbit_r48_c9 bl_9 br_9 wl_48 vdd gnd cell_6t
Xbit_r49_c9 bl_9 br_9 wl_49 vdd gnd cell_6t
Xbit_r50_c9 bl_9 br_9 wl_50 vdd gnd cell_6t
Xbit_r51_c9 bl_9 br_9 wl_51 vdd gnd cell_6t
Xbit_r52_c9 bl_9 br_9 wl_52 vdd gnd cell_6t
Xbit_r53_c9 bl_9 br_9 wl_53 vdd gnd cell_6t
Xbit_r54_c9 bl_9 br_9 wl_54 vdd gnd cell_6t
Xbit_r55_c9 bl_9 br_9 wl_55 vdd gnd cell_6t
Xbit_r56_c9 bl_9 br_9 wl_56 vdd gnd cell_6t
Xbit_r57_c9 bl_9 br_9 wl_57 vdd gnd cell_6t
Xbit_r58_c9 bl_9 br_9 wl_58 vdd gnd cell_6t
Xbit_r59_c9 bl_9 br_9 wl_59 vdd gnd cell_6t
Xbit_r60_c9 bl_9 br_9 wl_60 vdd gnd cell_6t
Xbit_r61_c9 bl_9 br_9 wl_61 vdd gnd cell_6t
Xbit_r62_c9 bl_9 br_9 wl_62 vdd gnd cell_6t
Xbit_r63_c9 bl_9 br_9 wl_63 vdd gnd cell_6t
Xbit_r64_c9 bl_9 br_9 wl_64 vdd gnd cell_6t
Xbit_r65_c9 bl_9 br_9 wl_65 vdd gnd cell_6t
Xbit_r66_c9 bl_9 br_9 wl_66 vdd gnd cell_6t
Xbit_r67_c9 bl_9 br_9 wl_67 vdd gnd cell_6t
Xbit_r68_c9 bl_9 br_9 wl_68 vdd gnd cell_6t
Xbit_r69_c9 bl_9 br_9 wl_69 vdd gnd cell_6t
Xbit_r70_c9 bl_9 br_9 wl_70 vdd gnd cell_6t
Xbit_r71_c9 bl_9 br_9 wl_71 vdd gnd cell_6t
Xbit_r72_c9 bl_9 br_9 wl_72 vdd gnd cell_6t
Xbit_r73_c9 bl_9 br_9 wl_73 vdd gnd cell_6t
Xbit_r74_c9 bl_9 br_9 wl_74 vdd gnd cell_6t
Xbit_r75_c9 bl_9 br_9 wl_75 vdd gnd cell_6t
Xbit_r76_c9 bl_9 br_9 wl_76 vdd gnd cell_6t
Xbit_r77_c9 bl_9 br_9 wl_77 vdd gnd cell_6t
Xbit_r78_c9 bl_9 br_9 wl_78 vdd gnd cell_6t
Xbit_r79_c9 bl_9 br_9 wl_79 vdd gnd cell_6t
Xbit_r80_c9 bl_9 br_9 wl_80 vdd gnd cell_6t
Xbit_r81_c9 bl_9 br_9 wl_81 vdd gnd cell_6t
Xbit_r82_c9 bl_9 br_9 wl_82 vdd gnd cell_6t
Xbit_r83_c9 bl_9 br_9 wl_83 vdd gnd cell_6t
Xbit_r84_c9 bl_9 br_9 wl_84 vdd gnd cell_6t
Xbit_r85_c9 bl_9 br_9 wl_85 vdd gnd cell_6t
Xbit_r86_c9 bl_9 br_9 wl_86 vdd gnd cell_6t
Xbit_r87_c9 bl_9 br_9 wl_87 vdd gnd cell_6t
Xbit_r88_c9 bl_9 br_9 wl_88 vdd gnd cell_6t
Xbit_r89_c9 bl_9 br_9 wl_89 vdd gnd cell_6t
Xbit_r90_c9 bl_9 br_9 wl_90 vdd gnd cell_6t
Xbit_r91_c9 bl_9 br_9 wl_91 vdd gnd cell_6t
Xbit_r92_c9 bl_9 br_9 wl_92 vdd gnd cell_6t
Xbit_r93_c9 bl_9 br_9 wl_93 vdd gnd cell_6t
Xbit_r94_c9 bl_9 br_9 wl_94 vdd gnd cell_6t
Xbit_r95_c9 bl_9 br_9 wl_95 vdd gnd cell_6t
Xbit_r96_c9 bl_9 br_9 wl_96 vdd gnd cell_6t
Xbit_r97_c9 bl_9 br_9 wl_97 vdd gnd cell_6t
Xbit_r98_c9 bl_9 br_9 wl_98 vdd gnd cell_6t
Xbit_r99_c9 bl_9 br_9 wl_99 vdd gnd cell_6t
Xbit_r100_c9 bl_9 br_9 wl_100 vdd gnd cell_6t
Xbit_r101_c9 bl_9 br_9 wl_101 vdd gnd cell_6t
Xbit_r102_c9 bl_9 br_9 wl_102 vdd gnd cell_6t
Xbit_r103_c9 bl_9 br_9 wl_103 vdd gnd cell_6t
Xbit_r104_c9 bl_9 br_9 wl_104 vdd gnd cell_6t
Xbit_r105_c9 bl_9 br_9 wl_105 vdd gnd cell_6t
Xbit_r106_c9 bl_9 br_9 wl_106 vdd gnd cell_6t
Xbit_r107_c9 bl_9 br_9 wl_107 vdd gnd cell_6t
Xbit_r108_c9 bl_9 br_9 wl_108 vdd gnd cell_6t
Xbit_r109_c9 bl_9 br_9 wl_109 vdd gnd cell_6t
Xbit_r110_c9 bl_9 br_9 wl_110 vdd gnd cell_6t
Xbit_r111_c9 bl_9 br_9 wl_111 vdd gnd cell_6t
Xbit_r112_c9 bl_9 br_9 wl_112 vdd gnd cell_6t
Xbit_r113_c9 bl_9 br_9 wl_113 vdd gnd cell_6t
Xbit_r114_c9 bl_9 br_9 wl_114 vdd gnd cell_6t
Xbit_r115_c9 bl_9 br_9 wl_115 vdd gnd cell_6t
Xbit_r116_c9 bl_9 br_9 wl_116 vdd gnd cell_6t
Xbit_r117_c9 bl_9 br_9 wl_117 vdd gnd cell_6t
Xbit_r118_c9 bl_9 br_9 wl_118 vdd gnd cell_6t
Xbit_r119_c9 bl_9 br_9 wl_119 vdd gnd cell_6t
Xbit_r120_c9 bl_9 br_9 wl_120 vdd gnd cell_6t
Xbit_r121_c9 bl_9 br_9 wl_121 vdd gnd cell_6t
Xbit_r122_c9 bl_9 br_9 wl_122 vdd gnd cell_6t
Xbit_r123_c9 bl_9 br_9 wl_123 vdd gnd cell_6t
Xbit_r124_c9 bl_9 br_9 wl_124 vdd gnd cell_6t
Xbit_r125_c9 bl_9 br_9 wl_125 vdd gnd cell_6t
Xbit_r126_c9 bl_9 br_9 wl_126 vdd gnd cell_6t
Xbit_r127_c9 bl_9 br_9 wl_127 vdd gnd cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd cell_6t
Xbit_r1_c10 bl_10 br_10 wl_1 vdd gnd cell_6t
Xbit_r2_c10 bl_10 br_10 wl_2 vdd gnd cell_6t
Xbit_r3_c10 bl_10 br_10 wl_3 vdd gnd cell_6t
Xbit_r4_c10 bl_10 br_10 wl_4 vdd gnd cell_6t
Xbit_r5_c10 bl_10 br_10 wl_5 vdd gnd cell_6t
Xbit_r6_c10 bl_10 br_10 wl_6 vdd gnd cell_6t
Xbit_r7_c10 bl_10 br_10 wl_7 vdd gnd cell_6t
Xbit_r8_c10 bl_10 br_10 wl_8 vdd gnd cell_6t
Xbit_r9_c10 bl_10 br_10 wl_9 vdd gnd cell_6t
Xbit_r10_c10 bl_10 br_10 wl_10 vdd gnd cell_6t
Xbit_r11_c10 bl_10 br_10 wl_11 vdd gnd cell_6t
Xbit_r12_c10 bl_10 br_10 wl_12 vdd gnd cell_6t
Xbit_r13_c10 bl_10 br_10 wl_13 vdd gnd cell_6t
Xbit_r14_c10 bl_10 br_10 wl_14 vdd gnd cell_6t
Xbit_r15_c10 bl_10 br_10 wl_15 vdd gnd cell_6t
Xbit_r16_c10 bl_10 br_10 wl_16 vdd gnd cell_6t
Xbit_r17_c10 bl_10 br_10 wl_17 vdd gnd cell_6t
Xbit_r18_c10 bl_10 br_10 wl_18 vdd gnd cell_6t
Xbit_r19_c10 bl_10 br_10 wl_19 vdd gnd cell_6t
Xbit_r20_c10 bl_10 br_10 wl_20 vdd gnd cell_6t
Xbit_r21_c10 bl_10 br_10 wl_21 vdd gnd cell_6t
Xbit_r22_c10 bl_10 br_10 wl_22 vdd gnd cell_6t
Xbit_r23_c10 bl_10 br_10 wl_23 vdd gnd cell_6t
Xbit_r24_c10 bl_10 br_10 wl_24 vdd gnd cell_6t
Xbit_r25_c10 bl_10 br_10 wl_25 vdd gnd cell_6t
Xbit_r26_c10 bl_10 br_10 wl_26 vdd gnd cell_6t
Xbit_r27_c10 bl_10 br_10 wl_27 vdd gnd cell_6t
Xbit_r28_c10 bl_10 br_10 wl_28 vdd gnd cell_6t
Xbit_r29_c10 bl_10 br_10 wl_29 vdd gnd cell_6t
Xbit_r30_c10 bl_10 br_10 wl_30 vdd gnd cell_6t
Xbit_r31_c10 bl_10 br_10 wl_31 vdd gnd cell_6t
Xbit_r32_c10 bl_10 br_10 wl_32 vdd gnd cell_6t
Xbit_r33_c10 bl_10 br_10 wl_33 vdd gnd cell_6t
Xbit_r34_c10 bl_10 br_10 wl_34 vdd gnd cell_6t
Xbit_r35_c10 bl_10 br_10 wl_35 vdd gnd cell_6t
Xbit_r36_c10 bl_10 br_10 wl_36 vdd gnd cell_6t
Xbit_r37_c10 bl_10 br_10 wl_37 vdd gnd cell_6t
Xbit_r38_c10 bl_10 br_10 wl_38 vdd gnd cell_6t
Xbit_r39_c10 bl_10 br_10 wl_39 vdd gnd cell_6t
Xbit_r40_c10 bl_10 br_10 wl_40 vdd gnd cell_6t
Xbit_r41_c10 bl_10 br_10 wl_41 vdd gnd cell_6t
Xbit_r42_c10 bl_10 br_10 wl_42 vdd gnd cell_6t
Xbit_r43_c10 bl_10 br_10 wl_43 vdd gnd cell_6t
Xbit_r44_c10 bl_10 br_10 wl_44 vdd gnd cell_6t
Xbit_r45_c10 bl_10 br_10 wl_45 vdd gnd cell_6t
Xbit_r46_c10 bl_10 br_10 wl_46 vdd gnd cell_6t
Xbit_r47_c10 bl_10 br_10 wl_47 vdd gnd cell_6t
Xbit_r48_c10 bl_10 br_10 wl_48 vdd gnd cell_6t
Xbit_r49_c10 bl_10 br_10 wl_49 vdd gnd cell_6t
Xbit_r50_c10 bl_10 br_10 wl_50 vdd gnd cell_6t
Xbit_r51_c10 bl_10 br_10 wl_51 vdd gnd cell_6t
Xbit_r52_c10 bl_10 br_10 wl_52 vdd gnd cell_6t
Xbit_r53_c10 bl_10 br_10 wl_53 vdd gnd cell_6t
Xbit_r54_c10 bl_10 br_10 wl_54 vdd gnd cell_6t
Xbit_r55_c10 bl_10 br_10 wl_55 vdd gnd cell_6t
Xbit_r56_c10 bl_10 br_10 wl_56 vdd gnd cell_6t
Xbit_r57_c10 bl_10 br_10 wl_57 vdd gnd cell_6t
Xbit_r58_c10 bl_10 br_10 wl_58 vdd gnd cell_6t
Xbit_r59_c10 bl_10 br_10 wl_59 vdd gnd cell_6t
Xbit_r60_c10 bl_10 br_10 wl_60 vdd gnd cell_6t
Xbit_r61_c10 bl_10 br_10 wl_61 vdd gnd cell_6t
Xbit_r62_c10 bl_10 br_10 wl_62 vdd gnd cell_6t
Xbit_r63_c10 bl_10 br_10 wl_63 vdd gnd cell_6t
Xbit_r64_c10 bl_10 br_10 wl_64 vdd gnd cell_6t
Xbit_r65_c10 bl_10 br_10 wl_65 vdd gnd cell_6t
Xbit_r66_c10 bl_10 br_10 wl_66 vdd gnd cell_6t
Xbit_r67_c10 bl_10 br_10 wl_67 vdd gnd cell_6t
Xbit_r68_c10 bl_10 br_10 wl_68 vdd gnd cell_6t
Xbit_r69_c10 bl_10 br_10 wl_69 vdd gnd cell_6t
Xbit_r70_c10 bl_10 br_10 wl_70 vdd gnd cell_6t
Xbit_r71_c10 bl_10 br_10 wl_71 vdd gnd cell_6t
Xbit_r72_c10 bl_10 br_10 wl_72 vdd gnd cell_6t
Xbit_r73_c10 bl_10 br_10 wl_73 vdd gnd cell_6t
Xbit_r74_c10 bl_10 br_10 wl_74 vdd gnd cell_6t
Xbit_r75_c10 bl_10 br_10 wl_75 vdd gnd cell_6t
Xbit_r76_c10 bl_10 br_10 wl_76 vdd gnd cell_6t
Xbit_r77_c10 bl_10 br_10 wl_77 vdd gnd cell_6t
Xbit_r78_c10 bl_10 br_10 wl_78 vdd gnd cell_6t
Xbit_r79_c10 bl_10 br_10 wl_79 vdd gnd cell_6t
Xbit_r80_c10 bl_10 br_10 wl_80 vdd gnd cell_6t
Xbit_r81_c10 bl_10 br_10 wl_81 vdd gnd cell_6t
Xbit_r82_c10 bl_10 br_10 wl_82 vdd gnd cell_6t
Xbit_r83_c10 bl_10 br_10 wl_83 vdd gnd cell_6t
Xbit_r84_c10 bl_10 br_10 wl_84 vdd gnd cell_6t
Xbit_r85_c10 bl_10 br_10 wl_85 vdd gnd cell_6t
Xbit_r86_c10 bl_10 br_10 wl_86 vdd gnd cell_6t
Xbit_r87_c10 bl_10 br_10 wl_87 vdd gnd cell_6t
Xbit_r88_c10 bl_10 br_10 wl_88 vdd gnd cell_6t
Xbit_r89_c10 bl_10 br_10 wl_89 vdd gnd cell_6t
Xbit_r90_c10 bl_10 br_10 wl_90 vdd gnd cell_6t
Xbit_r91_c10 bl_10 br_10 wl_91 vdd gnd cell_6t
Xbit_r92_c10 bl_10 br_10 wl_92 vdd gnd cell_6t
Xbit_r93_c10 bl_10 br_10 wl_93 vdd gnd cell_6t
Xbit_r94_c10 bl_10 br_10 wl_94 vdd gnd cell_6t
Xbit_r95_c10 bl_10 br_10 wl_95 vdd gnd cell_6t
Xbit_r96_c10 bl_10 br_10 wl_96 vdd gnd cell_6t
Xbit_r97_c10 bl_10 br_10 wl_97 vdd gnd cell_6t
Xbit_r98_c10 bl_10 br_10 wl_98 vdd gnd cell_6t
Xbit_r99_c10 bl_10 br_10 wl_99 vdd gnd cell_6t
Xbit_r100_c10 bl_10 br_10 wl_100 vdd gnd cell_6t
Xbit_r101_c10 bl_10 br_10 wl_101 vdd gnd cell_6t
Xbit_r102_c10 bl_10 br_10 wl_102 vdd gnd cell_6t
Xbit_r103_c10 bl_10 br_10 wl_103 vdd gnd cell_6t
Xbit_r104_c10 bl_10 br_10 wl_104 vdd gnd cell_6t
Xbit_r105_c10 bl_10 br_10 wl_105 vdd gnd cell_6t
Xbit_r106_c10 bl_10 br_10 wl_106 vdd gnd cell_6t
Xbit_r107_c10 bl_10 br_10 wl_107 vdd gnd cell_6t
Xbit_r108_c10 bl_10 br_10 wl_108 vdd gnd cell_6t
Xbit_r109_c10 bl_10 br_10 wl_109 vdd gnd cell_6t
Xbit_r110_c10 bl_10 br_10 wl_110 vdd gnd cell_6t
Xbit_r111_c10 bl_10 br_10 wl_111 vdd gnd cell_6t
Xbit_r112_c10 bl_10 br_10 wl_112 vdd gnd cell_6t
Xbit_r113_c10 bl_10 br_10 wl_113 vdd gnd cell_6t
Xbit_r114_c10 bl_10 br_10 wl_114 vdd gnd cell_6t
Xbit_r115_c10 bl_10 br_10 wl_115 vdd gnd cell_6t
Xbit_r116_c10 bl_10 br_10 wl_116 vdd gnd cell_6t
Xbit_r117_c10 bl_10 br_10 wl_117 vdd gnd cell_6t
Xbit_r118_c10 bl_10 br_10 wl_118 vdd gnd cell_6t
Xbit_r119_c10 bl_10 br_10 wl_119 vdd gnd cell_6t
Xbit_r120_c10 bl_10 br_10 wl_120 vdd gnd cell_6t
Xbit_r121_c10 bl_10 br_10 wl_121 vdd gnd cell_6t
Xbit_r122_c10 bl_10 br_10 wl_122 vdd gnd cell_6t
Xbit_r123_c10 bl_10 br_10 wl_123 vdd gnd cell_6t
Xbit_r124_c10 bl_10 br_10 wl_124 vdd gnd cell_6t
Xbit_r125_c10 bl_10 br_10 wl_125 vdd gnd cell_6t
Xbit_r126_c10 bl_10 br_10 wl_126 vdd gnd cell_6t
Xbit_r127_c10 bl_10 br_10 wl_127 vdd gnd cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd cell_6t
Xbit_r1_c11 bl_11 br_11 wl_1 vdd gnd cell_6t
Xbit_r2_c11 bl_11 br_11 wl_2 vdd gnd cell_6t
Xbit_r3_c11 bl_11 br_11 wl_3 vdd gnd cell_6t
Xbit_r4_c11 bl_11 br_11 wl_4 vdd gnd cell_6t
Xbit_r5_c11 bl_11 br_11 wl_5 vdd gnd cell_6t
Xbit_r6_c11 bl_11 br_11 wl_6 vdd gnd cell_6t
Xbit_r7_c11 bl_11 br_11 wl_7 vdd gnd cell_6t
Xbit_r8_c11 bl_11 br_11 wl_8 vdd gnd cell_6t
Xbit_r9_c11 bl_11 br_11 wl_9 vdd gnd cell_6t
Xbit_r10_c11 bl_11 br_11 wl_10 vdd gnd cell_6t
Xbit_r11_c11 bl_11 br_11 wl_11 vdd gnd cell_6t
Xbit_r12_c11 bl_11 br_11 wl_12 vdd gnd cell_6t
Xbit_r13_c11 bl_11 br_11 wl_13 vdd gnd cell_6t
Xbit_r14_c11 bl_11 br_11 wl_14 vdd gnd cell_6t
Xbit_r15_c11 bl_11 br_11 wl_15 vdd gnd cell_6t
Xbit_r16_c11 bl_11 br_11 wl_16 vdd gnd cell_6t
Xbit_r17_c11 bl_11 br_11 wl_17 vdd gnd cell_6t
Xbit_r18_c11 bl_11 br_11 wl_18 vdd gnd cell_6t
Xbit_r19_c11 bl_11 br_11 wl_19 vdd gnd cell_6t
Xbit_r20_c11 bl_11 br_11 wl_20 vdd gnd cell_6t
Xbit_r21_c11 bl_11 br_11 wl_21 vdd gnd cell_6t
Xbit_r22_c11 bl_11 br_11 wl_22 vdd gnd cell_6t
Xbit_r23_c11 bl_11 br_11 wl_23 vdd gnd cell_6t
Xbit_r24_c11 bl_11 br_11 wl_24 vdd gnd cell_6t
Xbit_r25_c11 bl_11 br_11 wl_25 vdd gnd cell_6t
Xbit_r26_c11 bl_11 br_11 wl_26 vdd gnd cell_6t
Xbit_r27_c11 bl_11 br_11 wl_27 vdd gnd cell_6t
Xbit_r28_c11 bl_11 br_11 wl_28 vdd gnd cell_6t
Xbit_r29_c11 bl_11 br_11 wl_29 vdd gnd cell_6t
Xbit_r30_c11 bl_11 br_11 wl_30 vdd gnd cell_6t
Xbit_r31_c11 bl_11 br_11 wl_31 vdd gnd cell_6t
Xbit_r32_c11 bl_11 br_11 wl_32 vdd gnd cell_6t
Xbit_r33_c11 bl_11 br_11 wl_33 vdd gnd cell_6t
Xbit_r34_c11 bl_11 br_11 wl_34 vdd gnd cell_6t
Xbit_r35_c11 bl_11 br_11 wl_35 vdd gnd cell_6t
Xbit_r36_c11 bl_11 br_11 wl_36 vdd gnd cell_6t
Xbit_r37_c11 bl_11 br_11 wl_37 vdd gnd cell_6t
Xbit_r38_c11 bl_11 br_11 wl_38 vdd gnd cell_6t
Xbit_r39_c11 bl_11 br_11 wl_39 vdd gnd cell_6t
Xbit_r40_c11 bl_11 br_11 wl_40 vdd gnd cell_6t
Xbit_r41_c11 bl_11 br_11 wl_41 vdd gnd cell_6t
Xbit_r42_c11 bl_11 br_11 wl_42 vdd gnd cell_6t
Xbit_r43_c11 bl_11 br_11 wl_43 vdd gnd cell_6t
Xbit_r44_c11 bl_11 br_11 wl_44 vdd gnd cell_6t
Xbit_r45_c11 bl_11 br_11 wl_45 vdd gnd cell_6t
Xbit_r46_c11 bl_11 br_11 wl_46 vdd gnd cell_6t
Xbit_r47_c11 bl_11 br_11 wl_47 vdd gnd cell_6t
Xbit_r48_c11 bl_11 br_11 wl_48 vdd gnd cell_6t
Xbit_r49_c11 bl_11 br_11 wl_49 vdd gnd cell_6t
Xbit_r50_c11 bl_11 br_11 wl_50 vdd gnd cell_6t
Xbit_r51_c11 bl_11 br_11 wl_51 vdd gnd cell_6t
Xbit_r52_c11 bl_11 br_11 wl_52 vdd gnd cell_6t
Xbit_r53_c11 bl_11 br_11 wl_53 vdd gnd cell_6t
Xbit_r54_c11 bl_11 br_11 wl_54 vdd gnd cell_6t
Xbit_r55_c11 bl_11 br_11 wl_55 vdd gnd cell_6t
Xbit_r56_c11 bl_11 br_11 wl_56 vdd gnd cell_6t
Xbit_r57_c11 bl_11 br_11 wl_57 vdd gnd cell_6t
Xbit_r58_c11 bl_11 br_11 wl_58 vdd gnd cell_6t
Xbit_r59_c11 bl_11 br_11 wl_59 vdd gnd cell_6t
Xbit_r60_c11 bl_11 br_11 wl_60 vdd gnd cell_6t
Xbit_r61_c11 bl_11 br_11 wl_61 vdd gnd cell_6t
Xbit_r62_c11 bl_11 br_11 wl_62 vdd gnd cell_6t
Xbit_r63_c11 bl_11 br_11 wl_63 vdd gnd cell_6t
Xbit_r64_c11 bl_11 br_11 wl_64 vdd gnd cell_6t
Xbit_r65_c11 bl_11 br_11 wl_65 vdd gnd cell_6t
Xbit_r66_c11 bl_11 br_11 wl_66 vdd gnd cell_6t
Xbit_r67_c11 bl_11 br_11 wl_67 vdd gnd cell_6t
Xbit_r68_c11 bl_11 br_11 wl_68 vdd gnd cell_6t
Xbit_r69_c11 bl_11 br_11 wl_69 vdd gnd cell_6t
Xbit_r70_c11 bl_11 br_11 wl_70 vdd gnd cell_6t
Xbit_r71_c11 bl_11 br_11 wl_71 vdd gnd cell_6t
Xbit_r72_c11 bl_11 br_11 wl_72 vdd gnd cell_6t
Xbit_r73_c11 bl_11 br_11 wl_73 vdd gnd cell_6t
Xbit_r74_c11 bl_11 br_11 wl_74 vdd gnd cell_6t
Xbit_r75_c11 bl_11 br_11 wl_75 vdd gnd cell_6t
Xbit_r76_c11 bl_11 br_11 wl_76 vdd gnd cell_6t
Xbit_r77_c11 bl_11 br_11 wl_77 vdd gnd cell_6t
Xbit_r78_c11 bl_11 br_11 wl_78 vdd gnd cell_6t
Xbit_r79_c11 bl_11 br_11 wl_79 vdd gnd cell_6t
Xbit_r80_c11 bl_11 br_11 wl_80 vdd gnd cell_6t
Xbit_r81_c11 bl_11 br_11 wl_81 vdd gnd cell_6t
Xbit_r82_c11 bl_11 br_11 wl_82 vdd gnd cell_6t
Xbit_r83_c11 bl_11 br_11 wl_83 vdd gnd cell_6t
Xbit_r84_c11 bl_11 br_11 wl_84 vdd gnd cell_6t
Xbit_r85_c11 bl_11 br_11 wl_85 vdd gnd cell_6t
Xbit_r86_c11 bl_11 br_11 wl_86 vdd gnd cell_6t
Xbit_r87_c11 bl_11 br_11 wl_87 vdd gnd cell_6t
Xbit_r88_c11 bl_11 br_11 wl_88 vdd gnd cell_6t
Xbit_r89_c11 bl_11 br_11 wl_89 vdd gnd cell_6t
Xbit_r90_c11 bl_11 br_11 wl_90 vdd gnd cell_6t
Xbit_r91_c11 bl_11 br_11 wl_91 vdd gnd cell_6t
Xbit_r92_c11 bl_11 br_11 wl_92 vdd gnd cell_6t
Xbit_r93_c11 bl_11 br_11 wl_93 vdd gnd cell_6t
Xbit_r94_c11 bl_11 br_11 wl_94 vdd gnd cell_6t
Xbit_r95_c11 bl_11 br_11 wl_95 vdd gnd cell_6t
Xbit_r96_c11 bl_11 br_11 wl_96 vdd gnd cell_6t
Xbit_r97_c11 bl_11 br_11 wl_97 vdd gnd cell_6t
Xbit_r98_c11 bl_11 br_11 wl_98 vdd gnd cell_6t
Xbit_r99_c11 bl_11 br_11 wl_99 vdd gnd cell_6t
Xbit_r100_c11 bl_11 br_11 wl_100 vdd gnd cell_6t
Xbit_r101_c11 bl_11 br_11 wl_101 vdd gnd cell_6t
Xbit_r102_c11 bl_11 br_11 wl_102 vdd gnd cell_6t
Xbit_r103_c11 bl_11 br_11 wl_103 vdd gnd cell_6t
Xbit_r104_c11 bl_11 br_11 wl_104 vdd gnd cell_6t
Xbit_r105_c11 bl_11 br_11 wl_105 vdd gnd cell_6t
Xbit_r106_c11 bl_11 br_11 wl_106 vdd gnd cell_6t
Xbit_r107_c11 bl_11 br_11 wl_107 vdd gnd cell_6t
Xbit_r108_c11 bl_11 br_11 wl_108 vdd gnd cell_6t
Xbit_r109_c11 bl_11 br_11 wl_109 vdd gnd cell_6t
Xbit_r110_c11 bl_11 br_11 wl_110 vdd gnd cell_6t
Xbit_r111_c11 bl_11 br_11 wl_111 vdd gnd cell_6t
Xbit_r112_c11 bl_11 br_11 wl_112 vdd gnd cell_6t
Xbit_r113_c11 bl_11 br_11 wl_113 vdd gnd cell_6t
Xbit_r114_c11 bl_11 br_11 wl_114 vdd gnd cell_6t
Xbit_r115_c11 bl_11 br_11 wl_115 vdd gnd cell_6t
Xbit_r116_c11 bl_11 br_11 wl_116 vdd gnd cell_6t
Xbit_r117_c11 bl_11 br_11 wl_117 vdd gnd cell_6t
Xbit_r118_c11 bl_11 br_11 wl_118 vdd gnd cell_6t
Xbit_r119_c11 bl_11 br_11 wl_119 vdd gnd cell_6t
Xbit_r120_c11 bl_11 br_11 wl_120 vdd gnd cell_6t
Xbit_r121_c11 bl_11 br_11 wl_121 vdd gnd cell_6t
Xbit_r122_c11 bl_11 br_11 wl_122 vdd gnd cell_6t
Xbit_r123_c11 bl_11 br_11 wl_123 vdd gnd cell_6t
Xbit_r124_c11 bl_11 br_11 wl_124 vdd gnd cell_6t
Xbit_r125_c11 bl_11 br_11 wl_125 vdd gnd cell_6t
Xbit_r126_c11 bl_11 br_11 wl_126 vdd gnd cell_6t
Xbit_r127_c11 bl_11 br_11 wl_127 vdd gnd cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd cell_6t
Xbit_r1_c12 bl_12 br_12 wl_1 vdd gnd cell_6t
Xbit_r2_c12 bl_12 br_12 wl_2 vdd gnd cell_6t
Xbit_r3_c12 bl_12 br_12 wl_3 vdd gnd cell_6t
Xbit_r4_c12 bl_12 br_12 wl_4 vdd gnd cell_6t
Xbit_r5_c12 bl_12 br_12 wl_5 vdd gnd cell_6t
Xbit_r6_c12 bl_12 br_12 wl_6 vdd gnd cell_6t
Xbit_r7_c12 bl_12 br_12 wl_7 vdd gnd cell_6t
Xbit_r8_c12 bl_12 br_12 wl_8 vdd gnd cell_6t
Xbit_r9_c12 bl_12 br_12 wl_9 vdd gnd cell_6t
Xbit_r10_c12 bl_12 br_12 wl_10 vdd gnd cell_6t
Xbit_r11_c12 bl_12 br_12 wl_11 vdd gnd cell_6t
Xbit_r12_c12 bl_12 br_12 wl_12 vdd gnd cell_6t
Xbit_r13_c12 bl_12 br_12 wl_13 vdd gnd cell_6t
Xbit_r14_c12 bl_12 br_12 wl_14 vdd gnd cell_6t
Xbit_r15_c12 bl_12 br_12 wl_15 vdd gnd cell_6t
Xbit_r16_c12 bl_12 br_12 wl_16 vdd gnd cell_6t
Xbit_r17_c12 bl_12 br_12 wl_17 vdd gnd cell_6t
Xbit_r18_c12 bl_12 br_12 wl_18 vdd gnd cell_6t
Xbit_r19_c12 bl_12 br_12 wl_19 vdd gnd cell_6t
Xbit_r20_c12 bl_12 br_12 wl_20 vdd gnd cell_6t
Xbit_r21_c12 bl_12 br_12 wl_21 vdd gnd cell_6t
Xbit_r22_c12 bl_12 br_12 wl_22 vdd gnd cell_6t
Xbit_r23_c12 bl_12 br_12 wl_23 vdd gnd cell_6t
Xbit_r24_c12 bl_12 br_12 wl_24 vdd gnd cell_6t
Xbit_r25_c12 bl_12 br_12 wl_25 vdd gnd cell_6t
Xbit_r26_c12 bl_12 br_12 wl_26 vdd gnd cell_6t
Xbit_r27_c12 bl_12 br_12 wl_27 vdd gnd cell_6t
Xbit_r28_c12 bl_12 br_12 wl_28 vdd gnd cell_6t
Xbit_r29_c12 bl_12 br_12 wl_29 vdd gnd cell_6t
Xbit_r30_c12 bl_12 br_12 wl_30 vdd gnd cell_6t
Xbit_r31_c12 bl_12 br_12 wl_31 vdd gnd cell_6t
Xbit_r32_c12 bl_12 br_12 wl_32 vdd gnd cell_6t
Xbit_r33_c12 bl_12 br_12 wl_33 vdd gnd cell_6t
Xbit_r34_c12 bl_12 br_12 wl_34 vdd gnd cell_6t
Xbit_r35_c12 bl_12 br_12 wl_35 vdd gnd cell_6t
Xbit_r36_c12 bl_12 br_12 wl_36 vdd gnd cell_6t
Xbit_r37_c12 bl_12 br_12 wl_37 vdd gnd cell_6t
Xbit_r38_c12 bl_12 br_12 wl_38 vdd gnd cell_6t
Xbit_r39_c12 bl_12 br_12 wl_39 vdd gnd cell_6t
Xbit_r40_c12 bl_12 br_12 wl_40 vdd gnd cell_6t
Xbit_r41_c12 bl_12 br_12 wl_41 vdd gnd cell_6t
Xbit_r42_c12 bl_12 br_12 wl_42 vdd gnd cell_6t
Xbit_r43_c12 bl_12 br_12 wl_43 vdd gnd cell_6t
Xbit_r44_c12 bl_12 br_12 wl_44 vdd gnd cell_6t
Xbit_r45_c12 bl_12 br_12 wl_45 vdd gnd cell_6t
Xbit_r46_c12 bl_12 br_12 wl_46 vdd gnd cell_6t
Xbit_r47_c12 bl_12 br_12 wl_47 vdd gnd cell_6t
Xbit_r48_c12 bl_12 br_12 wl_48 vdd gnd cell_6t
Xbit_r49_c12 bl_12 br_12 wl_49 vdd gnd cell_6t
Xbit_r50_c12 bl_12 br_12 wl_50 vdd gnd cell_6t
Xbit_r51_c12 bl_12 br_12 wl_51 vdd gnd cell_6t
Xbit_r52_c12 bl_12 br_12 wl_52 vdd gnd cell_6t
Xbit_r53_c12 bl_12 br_12 wl_53 vdd gnd cell_6t
Xbit_r54_c12 bl_12 br_12 wl_54 vdd gnd cell_6t
Xbit_r55_c12 bl_12 br_12 wl_55 vdd gnd cell_6t
Xbit_r56_c12 bl_12 br_12 wl_56 vdd gnd cell_6t
Xbit_r57_c12 bl_12 br_12 wl_57 vdd gnd cell_6t
Xbit_r58_c12 bl_12 br_12 wl_58 vdd gnd cell_6t
Xbit_r59_c12 bl_12 br_12 wl_59 vdd gnd cell_6t
Xbit_r60_c12 bl_12 br_12 wl_60 vdd gnd cell_6t
Xbit_r61_c12 bl_12 br_12 wl_61 vdd gnd cell_6t
Xbit_r62_c12 bl_12 br_12 wl_62 vdd gnd cell_6t
Xbit_r63_c12 bl_12 br_12 wl_63 vdd gnd cell_6t
Xbit_r64_c12 bl_12 br_12 wl_64 vdd gnd cell_6t
Xbit_r65_c12 bl_12 br_12 wl_65 vdd gnd cell_6t
Xbit_r66_c12 bl_12 br_12 wl_66 vdd gnd cell_6t
Xbit_r67_c12 bl_12 br_12 wl_67 vdd gnd cell_6t
Xbit_r68_c12 bl_12 br_12 wl_68 vdd gnd cell_6t
Xbit_r69_c12 bl_12 br_12 wl_69 vdd gnd cell_6t
Xbit_r70_c12 bl_12 br_12 wl_70 vdd gnd cell_6t
Xbit_r71_c12 bl_12 br_12 wl_71 vdd gnd cell_6t
Xbit_r72_c12 bl_12 br_12 wl_72 vdd gnd cell_6t
Xbit_r73_c12 bl_12 br_12 wl_73 vdd gnd cell_6t
Xbit_r74_c12 bl_12 br_12 wl_74 vdd gnd cell_6t
Xbit_r75_c12 bl_12 br_12 wl_75 vdd gnd cell_6t
Xbit_r76_c12 bl_12 br_12 wl_76 vdd gnd cell_6t
Xbit_r77_c12 bl_12 br_12 wl_77 vdd gnd cell_6t
Xbit_r78_c12 bl_12 br_12 wl_78 vdd gnd cell_6t
Xbit_r79_c12 bl_12 br_12 wl_79 vdd gnd cell_6t
Xbit_r80_c12 bl_12 br_12 wl_80 vdd gnd cell_6t
Xbit_r81_c12 bl_12 br_12 wl_81 vdd gnd cell_6t
Xbit_r82_c12 bl_12 br_12 wl_82 vdd gnd cell_6t
Xbit_r83_c12 bl_12 br_12 wl_83 vdd gnd cell_6t
Xbit_r84_c12 bl_12 br_12 wl_84 vdd gnd cell_6t
Xbit_r85_c12 bl_12 br_12 wl_85 vdd gnd cell_6t
Xbit_r86_c12 bl_12 br_12 wl_86 vdd gnd cell_6t
Xbit_r87_c12 bl_12 br_12 wl_87 vdd gnd cell_6t
Xbit_r88_c12 bl_12 br_12 wl_88 vdd gnd cell_6t
Xbit_r89_c12 bl_12 br_12 wl_89 vdd gnd cell_6t
Xbit_r90_c12 bl_12 br_12 wl_90 vdd gnd cell_6t
Xbit_r91_c12 bl_12 br_12 wl_91 vdd gnd cell_6t
Xbit_r92_c12 bl_12 br_12 wl_92 vdd gnd cell_6t
Xbit_r93_c12 bl_12 br_12 wl_93 vdd gnd cell_6t
Xbit_r94_c12 bl_12 br_12 wl_94 vdd gnd cell_6t
Xbit_r95_c12 bl_12 br_12 wl_95 vdd gnd cell_6t
Xbit_r96_c12 bl_12 br_12 wl_96 vdd gnd cell_6t
Xbit_r97_c12 bl_12 br_12 wl_97 vdd gnd cell_6t
Xbit_r98_c12 bl_12 br_12 wl_98 vdd gnd cell_6t
Xbit_r99_c12 bl_12 br_12 wl_99 vdd gnd cell_6t
Xbit_r100_c12 bl_12 br_12 wl_100 vdd gnd cell_6t
Xbit_r101_c12 bl_12 br_12 wl_101 vdd gnd cell_6t
Xbit_r102_c12 bl_12 br_12 wl_102 vdd gnd cell_6t
Xbit_r103_c12 bl_12 br_12 wl_103 vdd gnd cell_6t
Xbit_r104_c12 bl_12 br_12 wl_104 vdd gnd cell_6t
Xbit_r105_c12 bl_12 br_12 wl_105 vdd gnd cell_6t
Xbit_r106_c12 bl_12 br_12 wl_106 vdd gnd cell_6t
Xbit_r107_c12 bl_12 br_12 wl_107 vdd gnd cell_6t
Xbit_r108_c12 bl_12 br_12 wl_108 vdd gnd cell_6t
Xbit_r109_c12 bl_12 br_12 wl_109 vdd gnd cell_6t
Xbit_r110_c12 bl_12 br_12 wl_110 vdd gnd cell_6t
Xbit_r111_c12 bl_12 br_12 wl_111 vdd gnd cell_6t
Xbit_r112_c12 bl_12 br_12 wl_112 vdd gnd cell_6t
Xbit_r113_c12 bl_12 br_12 wl_113 vdd gnd cell_6t
Xbit_r114_c12 bl_12 br_12 wl_114 vdd gnd cell_6t
Xbit_r115_c12 bl_12 br_12 wl_115 vdd gnd cell_6t
Xbit_r116_c12 bl_12 br_12 wl_116 vdd gnd cell_6t
Xbit_r117_c12 bl_12 br_12 wl_117 vdd gnd cell_6t
Xbit_r118_c12 bl_12 br_12 wl_118 vdd gnd cell_6t
Xbit_r119_c12 bl_12 br_12 wl_119 vdd gnd cell_6t
Xbit_r120_c12 bl_12 br_12 wl_120 vdd gnd cell_6t
Xbit_r121_c12 bl_12 br_12 wl_121 vdd gnd cell_6t
Xbit_r122_c12 bl_12 br_12 wl_122 vdd gnd cell_6t
Xbit_r123_c12 bl_12 br_12 wl_123 vdd gnd cell_6t
Xbit_r124_c12 bl_12 br_12 wl_124 vdd gnd cell_6t
Xbit_r125_c12 bl_12 br_12 wl_125 vdd gnd cell_6t
Xbit_r126_c12 bl_12 br_12 wl_126 vdd gnd cell_6t
Xbit_r127_c12 bl_12 br_12 wl_127 vdd gnd cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd cell_6t
Xbit_r1_c13 bl_13 br_13 wl_1 vdd gnd cell_6t
Xbit_r2_c13 bl_13 br_13 wl_2 vdd gnd cell_6t
Xbit_r3_c13 bl_13 br_13 wl_3 vdd gnd cell_6t
Xbit_r4_c13 bl_13 br_13 wl_4 vdd gnd cell_6t
Xbit_r5_c13 bl_13 br_13 wl_5 vdd gnd cell_6t
Xbit_r6_c13 bl_13 br_13 wl_6 vdd gnd cell_6t
Xbit_r7_c13 bl_13 br_13 wl_7 vdd gnd cell_6t
Xbit_r8_c13 bl_13 br_13 wl_8 vdd gnd cell_6t
Xbit_r9_c13 bl_13 br_13 wl_9 vdd gnd cell_6t
Xbit_r10_c13 bl_13 br_13 wl_10 vdd gnd cell_6t
Xbit_r11_c13 bl_13 br_13 wl_11 vdd gnd cell_6t
Xbit_r12_c13 bl_13 br_13 wl_12 vdd gnd cell_6t
Xbit_r13_c13 bl_13 br_13 wl_13 vdd gnd cell_6t
Xbit_r14_c13 bl_13 br_13 wl_14 vdd gnd cell_6t
Xbit_r15_c13 bl_13 br_13 wl_15 vdd gnd cell_6t
Xbit_r16_c13 bl_13 br_13 wl_16 vdd gnd cell_6t
Xbit_r17_c13 bl_13 br_13 wl_17 vdd gnd cell_6t
Xbit_r18_c13 bl_13 br_13 wl_18 vdd gnd cell_6t
Xbit_r19_c13 bl_13 br_13 wl_19 vdd gnd cell_6t
Xbit_r20_c13 bl_13 br_13 wl_20 vdd gnd cell_6t
Xbit_r21_c13 bl_13 br_13 wl_21 vdd gnd cell_6t
Xbit_r22_c13 bl_13 br_13 wl_22 vdd gnd cell_6t
Xbit_r23_c13 bl_13 br_13 wl_23 vdd gnd cell_6t
Xbit_r24_c13 bl_13 br_13 wl_24 vdd gnd cell_6t
Xbit_r25_c13 bl_13 br_13 wl_25 vdd gnd cell_6t
Xbit_r26_c13 bl_13 br_13 wl_26 vdd gnd cell_6t
Xbit_r27_c13 bl_13 br_13 wl_27 vdd gnd cell_6t
Xbit_r28_c13 bl_13 br_13 wl_28 vdd gnd cell_6t
Xbit_r29_c13 bl_13 br_13 wl_29 vdd gnd cell_6t
Xbit_r30_c13 bl_13 br_13 wl_30 vdd gnd cell_6t
Xbit_r31_c13 bl_13 br_13 wl_31 vdd gnd cell_6t
Xbit_r32_c13 bl_13 br_13 wl_32 vdd gnd cell_6t
Xbit_r33_c13 bl_13 br_13 wl_33 vdd gnd cell_6t
Xbit_r34_c13 bl_13 br_13 wl_34 vdd gnd cell_6t
Xbit_r35_c13 bl_13 br_13 wl_35 vdd gnd cell_6t
Xbit_r36_c13 bl_13 br_13 wl_36 vdd gnd cell_6t
Xbit_r37_c13 bl_13 br_13 wl_37 vdd gnd cell_6t
Xbit_r38_c13 bl_13 br_13 wl_38 vdd gnd cell_6t
Xbit_r39_c13 bl_13 br_13 wl_39 vdd gnd cell_6t
Xbit_r40_c13 bl_13 br_13 wl_40 vdd gnd cell_6t
Xbit_r41_c13 bl_13 br_13 wl_41 vdd gnd cell_6t
Xbit_r42_c13 bl_13 br_13 wl_42 vdd gnd cell_6t
Xbit_r43_c13 bl_13 br_13 wl_43 vdd gnd cell_6t
Xbit_r44_c13 bl_13 br_13 wl_44 vdd gnd cell_6t
Xbit_r45_c13 bl_13 br_13 wl_45 vdd gnd cell_6t
Xbit_r46_c13 bl_13 br_13 wl_46 vdd gnd cell_6t
Xbit_r47_c13 bl_13 br_13 wl_47 vdd gnd cell_6t
Xbit_r48_c13 bl_13 br_13 wl_48 vdd gnd cell_6t
Xbit_r49_c13 bl_13 br_13 wl_49 vdd gnd cell_6t
Xbit_r50_c13 bl_13 br_13 wl_50 vdd gnd cell_6t
Xbit_r51_c13 bl_13 br_13 wl_51 vdd gnd cell_6t
Xbit_r52_c13 bl_13 br_13 wl_52 vdd gnd cell_6t
Xbit_r53_c13 bl_13 br_13 wl_53 vdd gnd cell_6t
Xbit_r54_c13 bl_13 br_13 wl_54 vdd gnd cell_6t
Xbit_r55_c13 bl_13 br_13 wl_55 vdd gnd cell_6t
Xbit_r56_c13 bl_13 br_13 wl_56 vdd gnd cell_6t
Xbit_r57_c13 bl_13 br_13 wl_57 vdd gnd cell_6t
Xbit_r58_c13 bl_13 br_13 wl_58 vdd gnd cell_6t
Xbit_r59_c13 bl_13 br_13 wl_59 vdd gnd cell_6t
Xbit_r60_c13 bl_13 br_13 wl_60 vdd gnd cell_6t
Xbit_r61_c13 bl_13 br_13 wl_61 vdd gnd cell_6t
Xbit_r62_c13 bl_13 br_13 wl_62 vdd gnd cell_6t
Xbit_r63_c13 bl_13 br_13 wl_63 vdd gnd cell_6t
Xbit_r64_c13 bl_13 br_13 wl_64 vdd gnd cell_6t
Xbit_r65_c13 bl_13 br_13 wl_65 vdd gnd cell_6t
Xbit_r66_c13 bl_13 br_13 wl_66 vdd gnd cell_6t
Xbit_r67_c13 bl_13 br_13 wl_67 vdd gnd cell_6t
Xbit_r68_c13 bl_13 br_13 wl_68 vdd gnd cell_6t
Xbit_r69_c13 bl_13 br_13 wl_69 vdd gnd cell_6t
Xbit_r70_c13 bl_13 br_13 wl_70 vdd gnd cell_6t
Xbit_r71_c13 bl_13 br_13 wl_71 vdd gnd cell_6t
Xbit_r72_c13 bl_13 br_13 wl_72 vdd gnd cell_6t
Xbit_r73_c13 bl_13 br_13 wl_73 vdd gnd cell_6t
Xbit_r74_c13 bl_13 br_13 wl_74 vdd gnd cell_6t
Xbit_r75_c13 bl_13 br_13 wl_75 vdd gnd cell_6t
Xbit_r76_c13 bl_13 br_13 wl_76 vdd gnd cell_6t
Xbit_r77_c13 bl_13 br_13 wl_77 vdd gnd cell_6t
Xbit_r78_c13 bl_13 br_13 wl_78 vdd gnd cell_6t
Xbit_r79_c13 bl_13 br_13 wl_79 vdd gnd cell_6t
Xbit_r80_c13 bl_13 br_13 wl_80 vdd gnd cell_6t
Xbit_r81_c13 bl_13 br_13 wl_81 vdd gnd cell_6t
Xbit_r82_c13 bl_13 br_13 wl_82 vdd gnd cell_6t
Xbit_r83_c13 bl_13 br_13 wl_83 vdd gnd cell_6t
Xbit_r84_c13 bl_13 br_13 wl_84 vdd gnd cell_6t
Xbit_r85_c13 bl_13 br_13 wl_85 vdd gnd cell_6t
Xbit_r86_c13 bl_13 br_13 wl_86 vdd gnd cell_6t
Xbit_r87_c13 bl_13 br_13 wl_87 vdd gnd cell_6t
Xbit_r88_c13 bl_13 br_13 wl_88 vdd gnd cell_6t
Xbit_r89_c13 bl_13 br_13 wl_89 vdd gnd cell_6t
Xbit_r90_c13 bl_13 br_13 wl_90 vdd gnd cell_6t
Xbit_r91_c13 bl_13 br_13 wl_91 vdd gnd cell_6t
Xbit_r92_c13 bl_13 br_13 wl_92 vdd gnd cell_6t
Xbit_r93_c13 bl_13 br_13 wl_93 vdd gnd cell_6t
Xbit_r94_c13 bl_13 br_13 wl_94 vdd gnd cell_6t
Xbit_r95_c13 bl_13 br_13 wl_95 vdd gnd cell_6t
Xbit_r96_c13 bl_13 br_13 wl_96 vdd gnd cell_6t
Xbit_r97_c13 bl_13 br_13 wl_97 vdd gnd cell_6t
Xbit_r98_c13 bl_13 br_13 wl_98 vdd gnd cell_6t
Xbit_r99_c13 bl_13 br_13 wl_99 vdd gnd cell_6t
Xbit_r100_c13 bl_13 br_13 wl_100 vdd gnd cell_6t
Xbit_r101_c13 bl_13 br_13 wl_101 vdd gnd cell_6t
Xbit_r102_c13 bl_13 br_13 wl_102 vdd gnd cell_6t
Xbit_r103_c13 bl_13 br_13 wl_103 vdd gnd cell_6t
Xbit_r104_c13 bl_13 br_13 wl_104 vdd gnd cell_6t
Xbit_r105_c13 bl_13 br_13 wl_105 vdd gnd cell_6t
Xbit_r106_c13 bl_13 br_13 wl_106 vdd gnd cell_6t
Xbit_r107_c13 bl_13 br_13 wl_107 vdd gnd cell_6t
Xbit_r108_c13 bl_13 br_13 wl_108 vdd gnd cell_6t
Xbit_r109_c13 bl_13 br_13 wl_109 vdd gnd cell_6t
Xbit_r110_c13 bl_13 br_13 wl_110 vdd gnd cell_6t
Xbit_r111_c13 bl_13 br_13 wl_111 vdd gnd cell_6t
Xbit_r112_c13 bl_13 br_13 wl_112 vdd gnd cell_6t
Xbit_r113_c13 bl_13 br_13 wl_113 vdd gnd cell_6t
Xbit_r114_c13 bl_13 br_13 wl_114 vdd gnd cell_6t
Xbit_r115_c13 bl_13 br_13 wl_115 vdd gnd cell_6t
Xbit_r116_c13 bl_13 br_13 wl_116 vdd gnd cell_6t
Xbit_r117_c13 bl_13 br_13 wl_117 vdd gnd cell_6t
Xbit_r118_c13 bl_13 br_13 wl_118 vdd gnd cell_6t
Xbit_r119_c13 bl_13 br_13 wl_119 vdd gnd cell_6t
Xbit_r120_c13 bl_13 br_13 wl_120 vdd gnd cell_6t
Xbit_r121_c13 bl_13 br_13 wl_121 vdd gnd cell_6t
Xbit_r122_c13 bl_13 br_13 wl_122 vdd gnd cell_6t
Xbit_r123_c13 bl_13 br_13 wl_123 vdd gnd cell_6t
Xbit_r124_c13 bl_13 br_13 wl_124 vdd gnd cell_6t
Xbit_r125_c13 bl_13 br_13 wl_125 vdd gnd cell_6t
Xbit_r126_c13 bl_13 br_13 wl_126 vdd gnd cell_6t
Xbit_r127_c13 bl_13 br_13 wl_127 vdd gnd cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd cell_6t
Xbit_r1_c14 bl_14 br_14 wl_1 vdd gnd cell_6t
Xbit_r2_c14 bl_14 br_14 wl_2 vdd gnd cell_6t
Xbit_r3_c14 bl_14 br_14 wl_3 vdd gnd cell_6t
Xbit_r4_c14 bl_14 br_14 wl_4 vdd gnd cell_6t
Xbit_r5_c14 bl_14 br_14 wl_5 vdd gnd cell_6t
Xbit_r6_c14 bl_14 br_14 wl_6 vdd gnd cell_6t
Xbit_r7_c14 bl_14 br_14 wl_7 vdd gnd cell_6t
Xbit_r8_c14 bl_14 br_14 wl_8 vdd gnd cell_6t
Xbit_r9_c14 bl_14 br_14 wl_9 vdd gnd cell_6t
Xbit_r10_c14 bl_14 br_14 wl_10 vdd gnd cell_6t
Xbit_r11_c14 bl_14 br_14 wl_11 vdd gnd cell_6t
Xbit_r12_c14 bl_14 br_14 wl_12 vdd gnd cell_6t
Xbit_r13_c14 bl_14 br_14 wl_13 vdd gnd cell_6t
Xbit_r14_c14 bl_14 br_14 wl_14 vdd gnd cell_6t
Xbit_r15_c14 bl_14 br_14 wl_15 vdd gnd cell_6t
Xbit_r16_c14 bl_14 br_14 wl_16 vdd gnd cell_6t
Xbit_r17_c14 bl_14 br_14 wl_17 vdd gnd cell_6t
Xbit_r18_c14 bl_14 br_14 wl_18 vdd gnd cell_6t
Xbit_r19_c14 bl_14 br_14 wl_19 vdd gnd cell_6t
Xbit_r20_c14 bl_14 br_14 wl_20 vdd gnd cell_6t
Xbit_r21_c14 bl_14 br_14 wl_21 vdd gnd cell_6t
Xbit_r22_c14 bl_14 br_14 wl_22 vdd gnd cell_6t
Xbit_r23_c14 bl_14 br_14 wl_23 vdd gnd cell_6t
Xbit_r24_c14 bl_14 br_14 wl_24 vdd gnd cell_6t
Xbit_r25_c14 bl_14 br_14 wl_25 vdd gnd cell_6t
Xbit_r26_c14 bl_14 br_14 wl_26 vdd gnd cell_6t
Xbit_r27_c14 bl_14 br_14 wl_27 vdd gnd cell_6t
Xbit_r28_c14 bl_14 br_14 wl_28 vdd gnd cell_6t
Xbit_r29_c14 bl_14 br_14 wl_29 vdd gnd cell_6t
Xbit_r30_c14 bl_14 br_14 wl_30 vdd gnd cell_6t
Xbit_r31_c14 bl_14 br_14 wl_31 vdd gnd cell_6t
Xbit_r32_c14 bl_14 br_14 wl_32 vdd gnd cell_6t
Xbit_r33_c14 bl_14 br_14 wl_33 vdd gnd cell_6t
Xbit_r34_c14 bl_14 br_14 wl_34 vdd gnd cell_6t
Xbit_r35_c14 bl_14 br_14 wl_35 vdd gnd cell_6t
Xbit_r36_c14 bl_14 br_14 wl_36 vdd gnd cell_6t
Xbit_r37_c14 bl_14 br_14 wl_37 vdd gnd cell_6t
Xbit_r38_c14 bl_14 br_14 wl_38 vdd gnd cell_6t
Xbit_r39_c14 bl_14 br_14 wl_39 vdd gnd cell_6t
Xbit_r40_c14 bl_14 br_14 wl_40 vdd gnd cell_6t
Xbit_r41_c14 bl_14 br_14 wl_41 vdd gnd cell_6t
Xbit_r42_c14 bl_14 br_14 wl_42 vdd gnd cell_6t
Xbit_r43_c14 bl_14 br_14 wl_43 vdd gnd cell_6t
Xbit_r44_c14 bl_14 br_14 wl_44 vdd gnd cell_6t
Xbit_r45_c14 bl_14 br_14 wl_45 vdd gnd cell_6t
Xbit_r46_c14 bl_14 br_14 wl_46 vdd gnd cell_6t
Xbit_r47_c14 bl_14 br_14 wl_47 vdd gnd cell_6t
Xbit_r48_c14 bl_14 br_14 wl_48 vdd gnd cell_6t
Xbit_r49_c14 bl_14 br_14 wl_49 vdd gnd cell_6t
Xbit_r50_c14 bl_14 br_14 wl_50 vdd gnd cell_6t
Xbit_r51_c14 bl_14 br_14 wl_51 vdd gnd cell_6t
Xbit_r52_c14 bl_14 br_14 wl_52 vdd gnd cell_6t
Xbit_r53_c14 bl_14 br_14 wl_53 vdd gnd cell_6t
Xbit_r54_c14 bl_14 br_14 wl_54 vdd gnd cell_6t
Xbit_r55_c14 bl_14 br_14 wl_55 vdd gnd cell_6t
Xbit_r56_c14 bl_14 br_14 wl_56 vdd gnd cell_6t
Xbit_r57_c14 bl_14 br_14 wl_57 vdd gnd cell_6t
Xbit_r58_c14 bl_14 br_14 wl_58 vdd gnd cell_6t
Xbit_r59_c14 bl_14 br_14 wl_59 vdd gnd cell_6t
Xbit_r60_c14 bl_14 br_14 wl_60 vdd gnd cell_6t
Xbit_r61_c14 bl_14 br_14 wl_61 vdd gnd cell_6t
Xbit_r62_c14 bl_14 br_14 wl_62 vdd gnd cell_6t
Xbit_r63_c14 bl_14 br_14 wl_63 vdd gnd cell_6t
Xbit_r64_c14 bl_14 br_14 wl_64 vdd gnd cell_6t
Xbit_r65_c14 bl_14 br_14 wl_65 vdd gnd cell_6t
Xbit_r66_c14 bl_14 br_14 wl_66 vdd gnd cell_6t
Xbit_r67_c14 bl_14 br_14 wl_67 vdd gnd cell_6t
Xbit_r68_c14 bl_14 br_14 wl_68 vdd gnd cell_6t
Xbit_r69_c14 bl_14 br_14 wl_69 vdd gnd cell_6t
Xbit_r70_c14 bl_14 br_14 wl_70 vdd gnd cell_6t
Xbit_r71_c14 bl_14 br_14 wl_71 vdd gnd cell_6t
Xbit_r72_c14 bl_14 br_14 wl_72 vdd gnd cell_6t
Xbit_r73_c14 bl_14 br_14 wl_73 vdd gnd cell_6t
Xbit_r74_c14 bl_14 br_14 wl_74 vdd gnd cell_6t
Xbit_r75_c14 bl_14 br_14 wl_75 vdd gnd cell_6t
Xbit_r76_c14 bl_14 br_14 wl_76 vdd gnd cell_6t
Xbit_r77_c14 bl_14 br_14 wl_77 vdd gnd cell_6t
Xbit_r78_c14 bl_14 br_14 wl_78 vdd gnd cell_6t
Xbit_r79_c14 bl_14 br_14 wl_79 vdd gnd cell_6t
Xbit_r80_c14 bl_14 br_14 wl_80 vdd gnd cell_6t
Xbit_r81_c14 bl_14 br_14 wl_81 vdd gnd cell_6t
Xbit_r82_c14 bl_14 br_14 wl_82 vdd gnd cell_6t
Xbit_r83_c14 bl_14 br_14 wl_83 vdd gnd cell_6t
Xbit_r84_c14 bl_14 br_14 wl_84 vdd gnd cell_6t
Xbit_r85_c14 bl_14 br_14 wl_85 vdd gnd cell_6t
Xbit_r86_c14 bl_14 br_14 wl_86 vdd gnd cell_6t
Xbit_r87_c14 bl_14 br_14 wl_87 vdd gnd cell_6t
Xbit_r88_c14 bl_14 br_14 wl_88 vdd gnd cell_6t
Xbit_r89_c14 bl_14 br_14 wl_89 vdd gnd cell_6t
Xbit_r90_c14 bl_14 br_14 wl_90 vdd gnd cell_6t
Xbit_r91_c14 bl_14 br_14 wl_91 vdd gnd cell_6t
Xbit_r92_c14 bl_14 br_14 wl_92 vdd gnd cell_6t
Xbit_r93_c14 bl_14 br_14 wl_93 vdd gnd cell_6t
Xbit_r94_c14 bl_14 br_14 wl_94 vdd gnd cell_6t
Xbit_r95_c14 bl_14 br_14 wl_95 vdd gnd cell_6t
Xbit_r96_c14 bl_14 br_14 wl_96 vdd gnd cell_6t
Xbit_r97_c14 bl_14 br_14 wl_97 vdd gnd cell_6t
Xbit_r98_c14 bl_14 br_14 wl_98 vdd gnd cell_6t
Xbit_r99_c14 bl_14 br_14 wl_99 vdd gnd cell_6t
Xbit_r100_c14 bl_14 br_14 wl_100 vdd gnd cell_6t
Xbit_r101_c14 bl_14 br_14 wl_101 vdd gnd cell_6t
Xbit_r102_c14 bl_14 br_14 wl_102 vdd gnd cell_6t
Xbit_r103_c14 bl_14 br_14 wl_103 vdd gnd cell_6t
Xbit_r104_c14 bl_14 br_14 wl_104 vdd gnd cell_6t
Xbit_r105_c14 bl_14 br_14 wl_105 vdd gnd cell_6t
Xbit_r106_c14 bl_14 br_14 wl_106 vdd gnd cell_6t
Xbit_r107_c14 bl_14 br_14 wl_107 vdd gnd cell_6t
Xbit_r108_c14 bl_14 br_14 wl_108 vdd gnd cell_6t
Xbit_r109_c14 bl_14 br_14 wl_109 vdd gnd cell_6t
Xbit_r110_c14 bl_14 br_14 wl_110 vdd gnd cell_6t
Xbit_r111_c14 bl_14 br_14 wl_111 vdd gnd cell_6t
Xbit_r112_c14 bl_14 br_14 wl_112 vdd gnd cell_6t
Xbit_r113_c14 bl_14 br_14 wl_113 vdd gnd cell_6t
Xbit_r114_c14 bl_14 br_14 wl_114 vdd gnd cell_6t
Xbit_r115_c14 bl_14 br_14 wl_115 vdd gnd cell_6t
Xbit_r116_c14 bl_14 br_14 wl_116 vdd gnd cell_6t
Xbit_r117_c14 bl_14 br_14 wl_117 vdd gnd cell_6t
Xbit_r118_c14 bl_14 br_14 wl_118 vdd gnd cell_6t
Xbit_r119_c14 bl_14 br_14 wl_119 vdd gnd cell_6t
Xbit_r120_c14 bl_14 br_14 wl_120 vdd gnd cell_6t
Xbit_r121_c14 bl_14 br_14 wl_121 vdd gnd cell_6t
Xbit_r122_c14 bl_14 br_14 wl_122 vdd gnd cell_6t
Xbit_r123_c14 bl_14 br_14 wl_123 vdd gnd cell_6t
Xbit_r124_c14 bl_14 br_14 wl_124 vdd gnd cell_6t
Xbit_r125_c14 bl_14 br_14 wl_125 vdd gnd cell_6t
Xbit_r126_c14 bl_14 br_14 wl_126 vdd gnd cell_6t
Xbit_r127_c14 bl_14 br_14 wl_127 vdd gnd cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd cell_6t
Xbit_r1_c15 bl_15 br_15 wl_1 vdd gnd cell_6t
Xbit_r2_c15 bl_15 br_15 wl_2 vdd gnd cell_6t
Xbit_r3_c15 bl_15 br_15 wl_3 vdd gnd cell_6t
Xbit_r4_c15 bl_15 br_15 wl_4 vdd gnd cell_6t
Xbit_r5_c15 bl_15 br_15 wl_5 vdd gnd cell_6t
Xbit_r6_c15 bl_15 br_15 wl_6 vdd gnd cell_6t
Xbit_r7_c15 bl_15 br_15 wl_7 vdd gnd cell_6t
Xbit_r8_c15 bl_15 br_15 wl_8 vdd gnd cell_6t
Xbit_r9_c15 bl_15 br_15 wl_9 vdd gnd cell_6t
Xbit_r10_c15 bl_15 br_15 wl_10 vdd gnd cell_6t
Xbit_r11_c15 bl_15 br_15 wl_11 vdd gnd cell_6t
Xbit_r12_c15 bl_15 br_15 wl_12 vdd gnd cell_6t
Xbit_r13_c15 bl_15 br_15 wl_13 vdd gnd cell_6t
Xbit_r14_c15 bl_15 br_15 wl_14 vdd gnd cell_6t
Xbit_r15_c15 bl_15 br_15 wl_15 vdd gnd cell_6t
Xbit_r16_c15 bl_15 br_15 wl_16 vdd gnd cell_6t
Xbit_r17_c15 bl_15 br_15 wl_17 vdd gnd cell_6t
Xbit_r18_c15 bl_15 br_15 wl_18 vdd gnd cell_6t
Xbit_r19_c15 bl_15 br_15 wl_19 vdd gnd cell_6t
Xbit_r20_c15 bl_15 br_15 wl_20 vdd gnd cell_6t
Xbit_r21_c15 bl_15 br_15 wl_21 vdd gnd cell_6t
Xbit_r22_c15 bl_15 br_15 wl_22 vdd gnd cell_6t
Xbit_r23_c15 bl_15 br_15 wl_23 vdd gnd cell_6t
Xbit_r24_c15 bl_15 br_15 wl_24 vdd gnd cell_6t
Xbit_r25_c15 bl_15 br_15 wl_25 vdd gnd cell_6t
Xbit_r26_c15 bl_15 br_15 wl_26 vdd gnd cell_6t
Xbit_r27_c15 bl_15 br_15 wl_27 vdd gnd cell_6t
Xbit_r28_c15 bl_15 br_15 wl_28 vdd gnd cell_6t
Xbit_r29_c15 bl_15 br_15 wl_29 vdd gnd cell_6t
Xbit_r30_c15 bl_15 br_15 wl_30 vdd gnd cell_6t
Xbit_r31_c15 bl_15 br_15 wl_31 vdd gnd cell_6t
Xbit_r32_c15 bl_15 br_15 wl_32 vdd gnd cell_6t
Xbit_r33_c15 bl_15 br_15 wl_33 vdd gnd cell_6t
Xbit_r34_c15 bl_15 br_15 wl_34 vdd gnd cell_6t
Xbit_r35_c15 bl_15 br_15 wl_35 vdd gnd cell_6t
Xbit_r36_c15 bl_15 br_15 wl_36 vdd gnd cell_6t
Xbit_r37_c15 bl_15 br_15 wl_37 vdd gnd cell_6t
Xbit_r38_c15 bl_15 br_15 wl_38 vdd gnd cell_6t
Xbit_r39_c15 bl_15 br_15 wl_39 vdd gnd cell_6t
Xbit_r40_c15 bl_15 br_15 wl_40 vdd gnd cell_6t
Xbit_r41_c15 bl_15 br_15 wl_41 vdd gnd cell_6t
Xbit_r42_c15 bl_15 br_15 wl_42 vdd gnd cell_6t
Xbit_r43_c15 bl_15 br_15 wl_43 vdd gnd cell_6t
Xbit_r44_c15 bl_15 br_15 wl_44 vdd gnd cell_6t
Xbit_r45_c15 bl_15 br_15 wl_45 vdd gnd cell_6t
Xbit_r46_c15 bl_15 br_15 wl_46 vdd gnd cell_6t
Xbit_r47_c15 bl_15 br_15 wl_47 vdd gnd cell_6t
Xbit_r48_c15 bl_15 br_15 wl_48 vdd gnd cell_6t
Xbit_r49_c15 bl_15 br_15 wl_49 vdd gnd cell_6t
Xbit_r50_c15 bl_15 br_15 wl_50 vdd gnd cell_6t
Xbit_r51_c15 bl_15 br_15 wl_51 vdd gnd cell_6t
Xbit_r52_c15 bl_15 br_15 wl_52 vdd gnd cell_6t
Xbit_r53_c15 bl_15 br_15 wl_53 vdd gnd cell_6t
Xbit_r54_c15 bl_15 br_15 wl_54 vdd gnd cell_6t
Xbit_r55_c15 bl_15 br_15 wl_55 vdd gnd cell_6t
Xbit_r56_c15 bl_15 br_15 wl_56 vdd gnd cell_6t
Xbit_r57_c15 bl_15 br_15 wl_57 vdd gnd cell_6t
Xbit_r58_c15 bl_15 br_15 wl_58 vdd gnd cell_6t
Xbit_r59_c15 bl_15 br_15 wl_59 vdd gnd cell_6t
Xbit_r60_c15 bl_15 br_15 wl_60 vdd gnd cell_6t
Xbit_r61_c15 bl_15 br_15 wl_61 vdd gnd cell_6t
Xbit_r62_c15 bl_15 br_15 wl_62 vdd gnd cell_6t
Xbit_r63_c15 bl_15 br_15 wl_63 vdd gnd cell_6t
Xbit_r64_c15 bl_15 br_15 wl_64 vdd gnd cell_6t
Xbit_r65_c15 bl_15 br_15 wl_65 vdd gnd cell_6t
Xbit_r66_c15 bl_15 br_15 wl_66 vdd gnd cell_6t
Xbit_r67_c15 bl_15 br_15 wl_67 vdd gnd cell_6t
Xbit_r68_c15 bl_15 br_15 wl_68 vdd gnd cell_6t
Xbit_r69_c15 bl_15 br_15 wl_69 vdd gnd cell_6t
Xbit_r70_c15 bl_15 br_15 wl_70 vdd gnd cell_6t
Xbit_r71_c15 bl_15 br_15 wl_71 vdd gnd cell_6t
Xbit_r72_c15 bl_15 br_15 wl_72 vdd gnd cell_6t
Xbit_r73_c15 bl_15 br_15 wl_73 vdd gnd cell_6t
Xbit_r74_c15 bl_15 br_15 wl_74 vdd gnd cell_6t
Xbit_r75_c15 bl_15 br_15 wl_75 vdd gnd cell_6t
Xbit_r76_c15 bl_15 br_15 wl_76 vdd gnd cell_6t
Xbit_r77_c15 bl_15 br_15 wl_77 vdd gnd cell_6t
Xbit_r78_c15 bl_15 br_15 wl_78 vdd gnd cell_6t
Xbit_r79_c15 bl_15 br_15 wl_79 vdd gnd cell_6t
Xbit_r80_c15 bl_15 br_15 wl_80 vdd gnd cell_6t
Xbit_r81_c15 bl_15 br_15 wl_81 vdd gnd cell_6t
Xbit_r82_c15 bl_15 br_15 wl_82 vdd gnd cell_6t
Xbit_r83_c15 bl_15 br_15 wl_83 vdd gnd cell_6t
Xbit_r84_c15 bl_15 br_15 wl_84 vdd gnd cell_6t
Xbit_r85_c15 bl_15 br_15 wl_85 vdd gnd cell_6t
Xbit_r86_c15 bl_15 br_15 wl_86 vdd gnd cell_6t
Xbit_r87_c15 bl_15 br_15 wl_87 vdd gnd cell_6t
Xbit_r88_c15 bl_15 br_15 wl_88 vdd gnd cell_6t
Xbit_r89_c15 bl_15 br_15 wl_89 vdd gnd cell_6t
Xbit_r90_c15 bl_15 br_15 wl_90 vdd gnd cell_6t
Xbit_r91_c15 bl_15 br_15 wl_91 vdd gnd cell_6t
Xbit_r92_c15 bl_15 br_15 wl_92 vdd gnd cell_6t
Xbit_r93_c15 bl_15 br_15 wl_93 vdd gnd cell_6t
Xbit_r94_c15 bl_15 br_15 wl_94 vdd gnd cell_6t
Xbit_r95_c15 bl_15 br_15 wl_95 vdd gnd cell_6t
Xbit_r96_c15 bl_15 br_15 wl_96 vdd gnd cell_6t
Xbit_r97_c15 bl_15 br_15 wl_97 vdd gnd cell_6t
Xbit_r98_c15 bl_15 br_15 wl_98 vdd gnd cell_6t
Xbit_r99_c15 bl_15 br_15 wl_99 vdd gnd cell_6t
Xbit_r100_c15 bl_15 br_15 wl_100 vdd gnd cell_6t
Xbit_r101_c15 bl_15 br_15 wl_101 vdd gnd cell_6t
Xbit_r102_c15 bl_15 br_15 wl_102 vdd gnd cell_6t
Xbit_r103_c15 bl_15 br_15 wl_103 vdd gnd cell_6t
Xbit_r104_c15 bl_15 br_15 wl_104 vdd gnd cell_6t
Xbit_r105_c15 bl_15 br_15 wl_105 vdd gnd cell_6t
Xbit_r106_c15 bl_15 br_15 wl_106 vdd gnd cell_6t
Xbit_r107_c15 bl_15 br_15 wl_107 vdd gnd cell_6t
Xbit_r108_c15 bl_15 br_15 wl_108 vdd gnd cell_6t
Xbit_r109_c15 bl_15 br_15 wl_109 vdd gnd cell_6t
Xbit_r110_c15 bl_15 br_15 wl_110 vdd gnd cell_6t
Xbit_r111_c15 bl_15 br_15 wl_111 vdd gnd cell_6t
Xbit_r112_c15 bl_15 br_15 wl_112 vdd gnd cell_6t
Xbit_r113_c15 bl_15 br_15 wl_113 vdd gnd cell_6t
Xbit_r114_c15 bl_15 br_15 wl_114 vdd gnd cell_6t
Xbit_r115_c15 bl_15 br_15 wl_115 vdd gnd cell_6t
Xbit_r116_c15 bl_15 br_15 wl_116 vdd gnd cell_6t
Xbit_r117_c15 bl_15 br_15 wl_117 vdd gnd cell_6t
Xbit_r118_c15 bl_15 br_15 wl_118 vdd gnd cell_6t
Xbit_r119_c15 bl_15 br_15 wl_119 vdd gnd cell_6t
Xbit_r120_c15 bl_15 br_15 wl_120 vdd gnd cell_6t
Xbit_r121_c15 bl_15 br_15 wl_121 vdd gnd cell_6t
Xbit_r122_c15 bl_15 br_15 wl_122 vdd gnd cell_6t
Xbit_r123_c15 bl_15 br_15 wl_123 vdd gnd cell_6t
Xbit_r124_c15 bl_15 br_15 wl_124 vdd gnd cell_6t
Xbit_r125_c15 bl_15 br_15 wl_125 vdd gnd cell_6t
Xbit_r126_c15 bl_15 br_15 wl_126 vdd gnd cell_6t
Xbit_r127_c15 bl_15 br_15 wl_127 vdd gnd cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd cell_6t
Xbit_r1_c16 bl_16 br_16 wl_1 vdd gnd cell_6t
Xbit_r2_c16 bl_16 br_16 wl_2 vdd gnd cell_6t
Xbit_r3_c16 bl_16 br_16 wl_3 vdd gnd cell_6t
Xbit_r4_c16 bl_16 br_16 wl_4 vdd gnd cell_6t
Xbit_r5_c16 bl_16 br_16 wl_5 vdd gnd cell_6t
Xbit_r6_c16 bl_16 br_16 wl_6 vdd gnd cell_6t
Xbit_r7_c16 bl_16 br_16 wl_7 vdd gnd cell_6t
Xbit_r8_c16 bl_16 br_16 wl_8 vdd gnd cell_6t
Xbit_r9_c16 bl_16 br_16 wl_9 vdd gnd cell_6t
Xbit_r10_c16 bl_16 br_16 wl_10 vdd gnd cell_6t
Xbit_r11_c16 bl_16 br_16 wl_11 vdd gnd cell_6t
Xbit_r12_c16 bl_16 br_16 wl_12 vdd gnd cell_6t
Xbit_r13_c16 bl_16 br_16 wl_13 vdd gnd cell_6t
Xbit_r14_c16 bl_16 br_16 wl_14 vdd gnd cell_6t
Xbit_r15_c16 bl_16 br_16 wl_15 vdd gnd cell_6t
Xbit_r16_c16 bl_16 br_16 wl_16 vdd gnd cell_6t
Xbit_r17_c16 bl_16 br_16 wl_17 vdd gnd cell_6t
Xbit_r18_c16 bl_16 br_16 wl_18 vdd gnd cell_6t
Xbit_r19_c16 bl_16 br_16 wl_19 vdd gnd cell_6t
Xbit_r20_c16 bl_16 br_16 wl_20 vdd gnd cell_6t
Xbit_r21_c16 bl_16 br_16 wl_21 vdd gnd cell_6t
Xbit_r22_c16 bl_16 br_16 wl_22 vdd gnd cell_6t
Xbit_r23_c16 bl_16 br_16 wl_23 vdd gnd cell_6t
Xbit_r24_c16 bl_16 br_16 wl_24 vdd gnd cell_6t
Xbit_r25_c16 bl_16 br_16 wl_25 vdd gnd cell_6t
Xbit_r26_c16 bl_16 br_16 wl_26 vdd gnd cell_6t
Xbit_r27_c16 bl_16 br_16 wl_27 vdd gnd cell_6t
Xbit_r28_c16 bl_16 br_16 wl_28 vdd gnd cell_6t
Xbit_r29_c16 bl_16 br_16 wl_29 vdd gnd cell_6t
Xbit_r30_c16 bl_16 br_16 wl_30 vdd gnd cell_6t
Xbit_r31_c16 bl_16 br_16 wl_31 vdd gnd cell_6t
Xbit_r32_c16 bl_16 br_16 wl_32 vdd gnd cell_6t
Xbit_r33_c16 bl_16 br_16 wl_33 vdd gnd cell_6t
Xbit_r34_c16 bl_16 br_16 wl_34 vdd gnd cell_6t
Xbit_r35_c16 bl_16 br_16 wl_35 vdd gnd cell_6t
Xbit_r36_c16 bl_16 br_16 wl_36 vdd gnd cell_6t
Xbit_r37_c16 bl_16 br_16 wl_37 vdd gnd cell_6t
Xbit_r38_c16 bl_16 br_16 wl_38 vdd gnd cell_6t
Xbit_r39_c16 bl_16 br_16 wl_39 vdd gnd cell_6t
Xbit_r40_c16 bl_16 br_16 wl_40 vdd gnd cell_6t
Xbit_r41_c16 bl_16 br_16 wl_41 vdd gnd cell_6t
Xbit_r42_c16 bl_16 br_16 wl_42 vdd gnd cell_6t
Xbit_r43_c16 bl_16 br_16 wl_43 vdd gnd cell_6t
Xbit_r44_c16 bl_16 br_16 wl_44 vdd gnd cell_6t
Xbit_r45_c16 bl_16 br_16 wl_45 vdd gnd cell_6t
Xbit_r46_c16 bl_16 br_16 wl_46 vdd gnd cell_6t
Xbit_r47_c16 bl_16 br_16 wl_47 vdd gnd cell_6t
Xbit_r48_c16 bl_16 br_16 wl_48 vdd gnd cell_6t
Xbit_r49_c16 bl_16 br_16 wl_49 vdd gnd cell_6t
Xbit_r50_c16 bl_16 br_16 wl_50 vdd gnd cell_6t
Xbit_r51_c16 bl_16 br_16 wl_51 vdd gnd cell_6t
Xbit_r52_c16 bl_16 br_16 wl_52 vdd gnd cell_6t
Xbit_r53_c16 bl_16 br_16 wl_53 vdd gnd cell_6t
Xbit_r54_c16 bl_16 br_16 wl_54 vdd gnd cell_6t
Xbit_r55_c16 bl_16 br_16 wl_55 vdd gnd cell_6t
Xbit_r56_c16 bl_16 br_16 wl_56 vdd gnd cell_6t
Xbit_r57_c16 bl_16 br_16 wl_57 vdd gnd cell_6t
Xbit_r58_c16 bl_16 br_16 wl_58 vdd gnd cell_6t
Xbit_r59_c16 bl_16 br_16 wl_59 vdd gnd cell_6t
Xbit_r60_c16 bl_16 br_16 wl_60 vdd gnd cell_6t
Xbit_r61_c16 bl_16 br_16 wl_61 vdd gnd cell_6t
Xbit_r62_c16 bl_16 br_16 wl_62 vdd gnd cell_6t
Xbit_r63_c16 bl_16 br_16 wl_63 vdd gnd cell_6t
Xbit_r64_c16 bl_16 br_16 wl_64 vdd gnd cell_6t
Xbit_r65_c16 bl_16 br_16 wl_65 vdd gnd cell_6t
Xbit_r66_c16 bl_16 br_16 wl_66 vdd gnd cell_6t
Xbit_r67_c16 bl_16 br_16 wl_67 vdd gnd cell_6t
Xbit_r68_c16 bl_16 br_16 wl_68 vdd gnd cell_6t
Xbit_r69_c16 bl_16 br_16 wl_69 vdd gnd cell_6t
Xbit_r70_c16 bl_16 br_16 wl_70 vdd gnd cell_6t
Xbit_r71_c16 bl_16 br_16 wl_71 vdd gnd cell_6t
Xbit_r72_c16 bl_16 br_16 wl_72 vdd gnd cell_6t
Xbit_r73_c16 bl_16 br_16 wl_73 vdd gnd cell_6t
Xbit_r74_c16 bl_16 br_16 wl_74 vdd gnd cell_6t
Xbit_r75_c16 bl_16 br_16 wl_75 vdd gnd cell_6t
Xbit_r76_c16 bl_16 br_16 wl_76 vdd gnd cell_6t
Xbit_r77_c16 bl_16 br_16 wl_77 vdd gnd cell_6t
Xbit_r78_c16 bl_16 br_16 wl_78 vdd gnd cell_6t
Xbit_r79_c16 bl_16 br_16 wl_79 vdd gnd cell_6t
Xbit_r80_c16 bl_16 br_16 wl_80 vdd gnd cell_6t
Xbit_r81_c16 bl_16 br_16 wl_81 vdd gnd cell_6t
Xbit_r82_c16 bl_16 br_16 wl_82 vdd gnd cell_6t
Xbit_r83_c16 bl_16 br_16 wl_83 vdd gnd cell_6t
Xbit_r84_c16 bl_16 br_16 wl_84 vdd gnd cell_6t
Xbit_r85_c16 bl_16 br_16 wl_85 vdd gnd cell_6t
Xbit_r86_c16 bl_16 br_16 wl_86 vdd gnd cell_6t
Xbit_r87_c16 bl_16 br_16 wl_87 vdd gnd cell_6t
Xbit_r88_c16 bl_16 br_16 wl_88 vdd gnd cell_6t
Xbit_r89_c16 bl_16 br_16 wl_89 vdd gnd cell_6t
Xbit_r90_c16 bl_16 br_16 wl_90 vdd gnd cell_6t
Xbit_r91_c16 bl_16 br_16 wl_91 vdd gnd cell_6t
Xbit_r92_c16 bl_16 br_16 wl_92 vdd gnd cell_6t
Xbit_r93_c16 bl_16 br_16 wl_93 vdd gnd cell_6t
Xbit_r94_c16 bl_16 br_16 wl_94 vdd gnd cell_6t
Xbit_r95_c16 bl_16 br_16 wl_95 vdd gnd cell_6t
Xbit_r96_c16 bl_16 br_16 wl_96 vdd gnd cell_6t
Xbit_r97_c16 bl_16 br_16 wl_97 vdd gnd cell_6t
Xbit_r98_c16 bl_16 br_16 wl_98 vdd gnd cell_6t
Xbit_r99_c16 bl_16 br_16 wl_99 vdd gnd cell_6t
Xbit_r100_c16 bl_16 br_16 wl_100 vdd gnd cell_6t
Xbit_r101_c16 bl_16 br_16 wl_101 vdd gnd cell_6t
Xbit_r102_c16 bl_16 br_16 wl_102 vdd gnd cell_6t
Xbit_r103_c16 bl_16 br_16 wl_103 vdd gnd cell_6t
Xbit_r104_c16 bl_16 br_16 wl_104 vdd gnd cell_6t
Xbit_r105_c16 bl_16 br_16 wl_105 vdd gnd cell_6t
Xbit_r106_c16 bl_16 br_16 wl_106 vdd gnd cell_6t
Xbit_r107_c16 bl_16 br_16 wl_107 vdd gnd cell_6t
Xbit_r108_c16 bl_16 br_16 wl_108 vdd gnd cell_6t
Xbit_r109_c16 bl_16 br_16 wl_109 vdd gnd cell_6t
Xbit_r110_c16 bl_16 br_16 wl_110 vdd gnd cell_6t
Xbit_r111_c16 bl_16 br_16 wl_111 vdd gnd cell_6t
Xbit_r112_c16 bl_16 br_16 wl_112 vdd gnd cell_6t
Xbit_r113_c16 bl_16 br_16 wl_113 vdd gnd cell_6t
Xbit_r114_c16 bl_16 br_16 wl_114 vdd gnd cell_6t
Xbit_r115_c16 bl_16 br_16 wl_115 vdd gnd cell_6t
Xbit_r116_c16 bl_16 br_16 wl_116 vdd gnd cell_6t
Xbit_r117_c16 bl_16 br_16 wl_117 vdd gnd cell_6t
Xbit_r118_c16 bl_16 br_16 wl_118 vdd gnd cell_6t
Xbit_r119_c16 bl_16 br_16 wl_119 vdd gnd cell_6t
Xbit_r120_c16 bl_16 br_16 wl_120 vdd gnd cell_6t
Xbit_r121_c16 bl_16 br_16 wl_121 vdd gnd cell_6t
Xbit_r122_c16 bl_16 br_16 wl_122 vdd gnd cell_6t
Xbit_r123_c16 bl_16 br_16 wl_123 vdd gnd cell_6t
Xbit_r124_c16 bl_16 br_16 wl_124 vdd gnd cell_6t
Xbit_r125_c16 bl_16 br_16 wl_125 vdd gnd cell_6t
Xbit_r126_c16 bl_16 br_16 wl_126 vdd gnd cell_6t
Xbit_r127_c16 bl_16 br_16 wl_127 vdd gnd cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd cell_6t
Xbit_r1_c17 bl_17 br_17 wl_1 vdd gnd cell_6t
Xbit_r2_c17 bl_17 br_17 wl_2 vdd gnd cell_6t
Xbit_r3_c17 bl_17 br_17 wl_3 vdd gnd cell_6t
Xbit_r4_c17 bl_17 br_17 wl_4 vdd gnd cell_6t
Xbit_r5_c17 bl_17 br_17 wl_5 vdd gnd cell_6t
Xbit_r6_c17 bl_17 br_17 wl_6 vdd gnd cell_6t
Xbit_r7_c17 bl_17 br_17 wl_7 vdd gnd cell_6t
Xbit_r8_c17 bl_17 br_17 wl_8 vdd gnd cell_6t
Xbit_r9_c17 bl_17 br_17 wl_9 vdd gnd cell_6t
Xbit_r10_c17 bl_17 br_17 wl_10 vdd gnd cell_6t
Xbit_r11_c17 bl_17 br_17 wl_11 vdd gnd cell_6t
Xbit_r12_c17 bl_17 br_17 wl_12 vdd gnd cell_6t
Xbit_r13_c17 bl_17 br_17 wl_13 vdd gnd cell_6t
Xbit_r14_c17 bl_17 br_17 wl_14 vdd gnd cell_6t
Xbit_r15_c17 bl_17 br_17 wl_15 vdd gnd cell_6t
Xbit_r16_c17 bl_17 br_17 wl_16 vdd gnd cell_6t
Xbit_r17_c17 bl_17 br_17 wl_17 vdd gnd cell_6t
Xbit_r18_c17 bl_17 br_17 wl_18 vdd gnd cell_6t
Xbit_r19_c17 bl_17 br_17 wl_19 vdd gnd cell_6t
Xbit_r20_c17 bl_17 br_17 wl_20 vdd gnd cell_6t
Xbit_r21_c17 bl_17 br_17 wl_21 vdd gnd cell_6t
Xbit_r22_c17 bl_17 br_17 wl_22 vdd gnd cell_6t
Xbit_r23_c17 bl_17 br_17 wl_23 vdd gnd cell_6t
Xbit_r24_c17 bl_17 br_17 wl_24 vdd gnd cell_6t
Xbit_r25_c17 bl_17 br_17 wl_25 vdd gnd cell_6t
Xbit_r26_c17 bl_17 br_17 wl_26 vdd gnd cell_6t
Xbit_r27_c17 bl_17 br_17 wl_27 vdd gnd cell_6t
Xbit_r28_c17 bl_17 br_17 wl_28 vdd gnd cell_6t
Xbit_r29_c17 bl_17 br_17 wl_29 vdd gnd cell_6t
Xbit_r30_c17 bl_17 br_17 wl_30 vdd gnd cell_6t
Xbit_r31_c17 bl_17 br_17 wl_31 vdd gnd cell_6t
Xbit_r32_c17 bl_17 br_17 wl_32 vdd gnd cell_6t
Xbit_r33_c17 bl_17 br_17 wl_33 vdd gnd cell_6t
Xbit_r34_c17 bl_17 br_17 wl_34 vdd gnd cell_6t
Xbit_r35_c17 bl_17 br_17 wl_35 vdd gnd cell_6t
Xbit_r36_c17 bl_17 br_17 wl_36 vdd gnd cell_6t
Xbit_r37_c17 bl_17 br_17 wl_37 vdd gnd cell_6t
Xbit_r38_c17 bl_17 br_17 wl_38 vdd gnd cell_6t
Xbit_r39_c17 bl_17 br_17 wl_39 vdd gnd cell_6t
Xbit_r40_c17 bl_17 br_17 wl_40 vdd gnd cell_6t
Xbit_r41_c17 bl_17 br_17 wl_41 vdd gnd cell_6t
Xbit_r42_c17 bl_17 br_17 wl_42 vdd gnd cell_6t
Xbit_r43_c17 bl_17 br_17 wl_43 vdd gnd cell_6t
Xbit_r44_c17 bl_17 br_17 wl_44 vdd gnd cell_6t
Xbit_r45_c17 bl_17 br_17 wl_45 vdd gnd cell_6t
Xbit_r46_c17 bl_17 br_17 wl_46 vdd gnd cell_6t
Xbit_r47_c17 bl_17 br_17 wl_47 vdd gnd cell_6t
Xbit_r48_c17 bl_17 br_17 wl_48 vdd gnd cell_6t
Xbit_r49_c17 bl_17 br_17 wl_49 vdd gnd cell_6t
Xbit_r50_c17 bl_17 br_17 wl_50 vdd gnd cell_6t
Xbit_r51_c17 bl_17 br_17 wl_51 vdd gnd cell_6t
Xbit_r52_c17 bl_17 br_17 wl_52 vdd gnd cell_6t
Xbit_r53_c17 bl_17 br_17 wl_53 vdd gnd cell_6t
Xbit_r54_c17 bl_17 br_17 wl_54 vdd gnd cell_6t
Xbit_r55_c17 bl_17 br_17 wl_55 vdd gnd cell_6t
Xbit_r56_c17 bl_17 br_17 wl_56 vdd gnd cell_6t
Xbit_r57_c17 bl_17 br_17 wl_57 vdd gnd cell_6t
Xbit_r58_c17 bl_17 br_17 wl_58 vdd gnd cell_6t
Xbit_r59_c17 bl_17 br_17 wl_59 vdd gnd cell_6t
Xbit_r60_c17 bl_17 br_17 wl_60 vdd gnd cell_6t
Xbit_r61_c17 bl_17 br_17 wl_61 vdd gnd cell_6t
Xbit_r62_c17 bl_17 br_17 wl_62 vdd gnd cell_6t
Xbit_r63_c17 bl_17 br_17 wl_63 vdd gnd cell_6t
Xbit_r64_c17 bl_17 br_17 wl_64 vdd gnd cell_6t
Xbit_r65_c17 bl_17 br_17 wl_65 vdd gnd cell_6t
Xbit_r66_c17 bl_17 br_17 wl_66 vdd gnd cell_6t
Xbit_r67_c17 bl_17 br_17 wl_67 vdd gnd cell_6t
Xbit_r68_c17 bl_17 br_17 wl_68 vdd gnd cell_6t
Xbit_r69_c17 bl_17 br_17 wl_69 vdd gnd cell_6t
Xbit_r70_c17 bl_17 br_17 wl_70 vdd gnd cell_6t
Xbit_r71_c17 bl_17 br_17 wl_71 vdd gnd cell_6t
Xbit_r72_c17 bl_17 br_17 wl_72 vdd gnd cell_6t
Xbit_r73_c17 bl_17 br_17 wl_73 vdd gnd cell_6t
Xbit_r74_c17 bl_17 br_17 wl_74 vdd gnd cell_6t
Xbit_r75_c17 bl_17 br_17 wl_75 vdd gnd cell_6t
Xbit_r76_c17 bl_17 br_17 wl_76 vdd gnd cell_6t
Xbit_r77_c17 bl_17 br_17 wl_77 vdd gnd cell_6t
Xbit_r78_c17 bl_17 br_17 wl_78 vdd gnd cell_6t
Xbit_r79_c17 bl_17 br_17 wl_79 vdd gnd cell_6t
Xbit_r80_c17 bl_17 br_17 wl_80 vdd gnd cell_6t
Xbit_r81_c17 bl_17 br_17 wl_81 vdd gnd cell_6t
Xbit_r82_c17 bl_17 br_17 wl_82 vdd gnd cell_6t
Xbit_r83_c17 bl_17 br_17 wl_83 vdd gnd cell_6t
Xbit_r84_c17 bl_17 br_17 wl_84 vdd gnd cell_6t
Xbit_r85_c17 bl_17 br_17 wl_85 vdd gnd cell_6t
Xbit_r86_c17 bl_17 br_17 wl_86 vdd gnd cell_6t
Xbit_r87_c17 bl_17 br_17 wl_87 vdd gnd cell_6t
Xbit_r88_c17 bl_17 br_17 wl_88 vdd gnd cell_6t
Xbit_r89_c17 bl_17 br_17 wl_89 vdd gnd cell_6t
Xbit_r90_c17 bl_17 br_17 wl_90 vdd gnd cell_6t
Xbit_r91_c17 bl_17 br_17 wl_91 vdd gnd cell_6t
Xbit_r92_c17 bl_17 br_17 wl_92 vdd gnd cell_6t
Xbit_r93_c17 bl_17 br_17 wl_93 vdd gnd cell_6t
Xbit_r94_c17 bl_17 br_17 wl_94 vdd gnd cell_6t
Xbit_r95_c17 bl_17 br_17 wl_95 vdd gnd cell_6t
Xbit_r96_c17 bl_17 br_17 wl_96 vdd gnd cell_6t
Xbit_r97_c17 bl_17 br_17 wl_97 vdd gnd cell_6t
Xbit_r98_c17 bl_17 br_17 wl_98 vdd gnd cell_6t
Xbit_r99_c17 bl_17 br_17 wl_99 vdd gnd cell_6t
Xbit_r100_c17 bl_17 br_17 wl_100 vdd gnd cell_6t
Xbit_r101_c17 bl_17 br_17 wl_101 vdd gnd cell_6t
Xbit_r102_c17 bl_17 br_17 wl_102 vdd gnd cell_6t
Xbit_r103_c17 bl_17 br_17 wl_103 vdd gnd cell_6t
Xbit_r104_c17 bl_17 br_17 wl_104 vdd gnd cell_6t
Xbit_r105_c17 bl_17 br_17 wl_105 vdd gnd cell_6t
Xbit_r106_c17 bl_17 br_17 wl_106 vdd gnd cell_6t
Xbit_r107_c17 bl_17 br_17 wl_107 vdd gnd cell_6t
Xbit_r108_c17 bl_17 br_17 wl_108 vdd gnd cell_6t
Xbit_r109_c17 bl_17 br_17 wl_109 vdd gnd cell_6t
Xbit_r110_c17 bl_17 br_17 wl_110 vdd gnd cell_6t
Xbit_r111_c17 bl_17 br_17 wl_111 vdd gnd cell_6t
Xbit_r112_c17 bl_17 br_17 wl_112 vdd gnd cell_6t
Xbit_r113_c17 bl_17 br_17 wl_113 vdd gnd cell_6t
Xbit_r114_c17 bl_17 br_17 wl_114 vdd gnd cell_6t
Xbit_r115_c17 bl_17 br_17 wl_115 vdd gnd cell_6t
Xbit_r116_c17 bl_17 br_17 wl_116 vdd gnd cell_6t
Xbit_r117_c17 bl_17 br_17 wl_117 vdd gnd cell_6t
Xbit_r118_c17 bl_17 br_17 wl_118 vdd gnd cell_6t
Xbit_r119_c17 bl_17 br_17 wl_119 vdd gnd cell_6t
Xbit_r120_c17 bl_17 br_17 wl_120 vdd gnd cell_6t
Xbit_r121_c17 bl_17 br_17 wl_121 vdd gnd cell_6t
Xbit_r122_c17 bl_17 br_17 wl_122 vdd gnd cell_6t
Xbit_r123_c17 bl_17 br_17 wl_123 vdd gnd cell_6t
Xbit_r124_c17 bl_17 br_17 wl_124 vdd gnd cell_6t
Xbit_r125_c17 bl_17 br_17 wl_125 vdd gnd cell_6t
Xbit_r126_c17 bl_17 br_17 wl_126 vdd gnd cell_6t
Xbit_r127_c17 bl_17 br_17 wl_127 vdd gnd cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd cell_6t
Xbit_r1_c18 bl_18 br_18 wl_1 vdd gnd cell_6t
Xbit_r2_c18 bl_18 br_18 wl_2 vdd gnd cell_6t
Xbit_r3_c18 bl_18 br_18 wl_3 vdd gnd cell_6t
Xbit_r4_c18 bl_18 br_18 wl_4 vdd gnd cell_6t
Xbit_r5_c18 bl_18 br_18 wl_5 vdd gnd cell_6t
Xbit_r6_c18 bl_18 br_18 wl_6 vdd gnd cell_6t
Xbit_r7_c18 bl_18 br_18 wl_7 vdd gnd cell_6t
Xbit_r8_c18 bl_18 br_18 wl_8 vdd gnd cell_6t
Xbit_r9_c18 bl_18 br_18 wl_9 vdd gnd cell_6t
Xbit_r10_c18 bl_18 br_18 wl_10 vdd gnd cell_6t
Xbit_r11_c18 bl_18 br_18 wl_11 vdd gnd cell_6t
Xbit_r12_c18 bl_18 br_18 wl_12 vdd gnd cell_6t
Xbit_r13_c18 bl_18 br_18 wl_13 vdd gnd cell_6t
Xbit_r14_c18 bl_18 br_18 wl_14 vdd gnd cell_6t
Xbit_r15_c18 bl_18 br_18 wl_15 vdd gnd cell_6t
Xbit_r16_c18 bl_18 br_18 wl_16 vdd gnd cell_6t
Xbit_r17_c18 bl_18 br_18 wl_17 vdd gnd cell_6t
Xbit_r18_c18 bl_18 br_18 wl_18 vdd gnd cell_6t
Xbit_r19_c18 bl_18 br_18 wl_19 vdd gnd cell_6t
Xbit_r20_c18 bl_18 br_18 wl_20 vdd gnd cell_6t
Xbit_r21_c18 bl_18 br_18 wl_21 vdd gnd cell_6t
Xbit_r22_c18 bl_18 br_18 wl_22 vdd gnd cell_6t
Xbit_r23_c18 bl_18 br_18 wl_23 vdd gnd cell_6t
Xbit_r24_c18 bl_18 br_18 wl_24 vdd gnd cell_6t
Xbit_r25_c18 bl_18 br_18 wl_25 vdd gnd cell_6t
Xbit_r26_c18 bl_18 br_18 wl_26 vdd gnd cell_6t
Xbit_r27_c18 bl_18 br_18 wl_27 vdd gnd cell_6t
Xbit_r28_c18 bl_18 br_18 wl_28 vdd gnd cell_6t
Xbit_r29_c18 bl_18 br_18 wl_29 vdd gnd cell_6t
Xbit_r30_c18 bl_18 br_18 wl_30 vdd gnd cell_6t
Xbit_r31_c18 bl_18 br_18 wl_31 vdd gnd cell_6t
Xbit_r32_c18 bl_18 br_18 wl_32 vdd gnd cell_6t
Xbit_r33_c18 bl_18 br_18 wl_33 vdd gnd cell_6t
Xbit_r34_c18 bl_18 br_18 wl_34 vdd gnd cell_6t
Xbit_r35_c18 bl_18 br_18 wl_35 vdd gnd cell_6t
Xbit_r36_c18 bl_18 br_18 wl_36 vdd gnd cell_6t
Xbit_r37_c18 bl_18 br_18 wl_37 vdd gnd cell_6t
Xbit_r38_c18 bl_18 br_18 wl_38 vdd gnd cell_6t
Xbit_r39_c18 bl_18 br_18 wl_39 vdd gnd cell_6t
Xbit_r40_c18 bl_18 br_18 wl_40 vdd gnd cell_6t
Xbit_r41_c18 bl_18 br_18 wl_41 vdd gnd cell_6t
Xbit_r42_c18 bl_18 br_18 wl_42 vdd gnd cell_6t
Xbit_r43_c18 bl_18 br_18 wl_43 vdd gnd cell_6t
Xbit_r44_c18 bl_18 br_18 wl_44 vdd gnd cell_6t
Xbit_r45_c18 bl_18 br_18 wl_45 vdd gnd cell_6t
Xbit_r46_c18 bl_18 br_18 wl_46 vdd gnd cell_6t
Xbit_r47_c18 bl_18 br_18 wl_47 vdd gnd cell_6t
Xbit_r48_c18 bl_18 br_18 wl_48 vdd gnd cell_6t
Xbit_r49_c18 bl_18 br_18 wl_49 vdd gnd cell_6t
Xbit_r50_c18 bl_18 br_18 wl_50 vdd gnd cell_6t
Xbit_r51_c18 bl_18 br_18 wl_51 vdd gnd cell_6t
Xbit_r52_c18 bl_18 br_18 wl_52 vdd gnd cell_6t
Xbit_r53_c18 bl_18 br_18 wl_53 vdd gnd cell_6t
Xbit_r54_c18 bl_18 br_18 wl_54 vdd gnd cell_6t
Xbit_r55_c18 bl_18 br_18 wl_55 vdd gnd cell_6t
Xbit_r56_c18 bl_18 br_18 wl_56 vdd gnd cell_6t
Xbit_r57_c18 bl_18 br_18 wl_57 vdd gnd cell_6t
Xbit_r58_c18 bl_18 br_18 wl_58 vdd gnd cell_6t
Xbit_r59_c18 bl_18 br_18 wl_59 vdd gnd cell_6t
Xbit_r60_c18 bl_18 br_18 wl_60 vdd gnd cell_6t
Xbit_r61_c18 bl_18 br_18 wl_61 vdd gnd cell_6t
Xbit_r62_c18 bl_18 br_18 wl_62 vdd gnd cell_6t
Xbit_r63_c18 bl_18 br_18 wl_63 vdd gnd cell_6t
Xbit_r64_c18 bl_18 br_18 wl_64 vdd gnd cell_6t
Xbit_r65_c18 bl_18 br_18 wl_65 vdd gnd cell_6t
Xbit_r66_c18 bl_18 br_18 wl_66 vdd gnd cell_6t
Xbit_r67_c18 bl_18 br_18 wl_67 vdd gnd cell_6t
Xbit_r68_c18 bl_18 br_18 wl_68 vdd gnd cell_6t
Xbit_r69_c18 bl_18 br_18 wl_69 vdd gnd cell_6t
Xbit_r70_c18 bl_18 br_18 wl_70 vdd gnd cell_6t
Xbit_r71_c18 bl_18 br_18 wl_71 vdd gnd cell_6t
Xbit_r72_c18 bl_18 br_18 wl_72 vdd gnd cell_6t
Xbit_r73_c18 bl_18 br_18 wl_73 vdd gnd cell_6t
Xbit_r74_c18 bl_18 br_18 wl_74 vdd gnd cell_6t
Xbit_r75_c18 bl_18 br_18 wl_75 vdd gnd cell_6t
Xbit_r76_c18 bl_18 br_18 wl_76 vdd gnd cell_6t
Xbit_r77_c18 bl_18 br_18 wl_77 vdd gnd cell_6t
Xbit_r78_c18 bl_18 br_18 wl_78 vdd gnd cell_6t
Xbit_r79_c18 bl_18 br_18 wl_79 vdd gnd cell_6t
Xbit_r80_c18 bl_18 br_18 wl_80 vdd gnd cell_6t
Xbit_r81_c18 bl_18 br_18 wl_81 vdd gnd cell_6t
Xbit_r82_c18 bl_18 br_18 wl_82 vdd gnd cell_6t
Xbit_r83_c18 bl_18 br_18 wl_83 vdd gnd cell_6t
Xbit_r84_c18 bl_18 br_18 wl_84 vdd gnd cell_6t
Xbit_r85_c18 bl_18 br_18 wl_85 vdd gnd cell_6t
Xbit_r86_c18 bl_18 br_18 wl_86 vdd gnd cell_6t
Xbit_r87_c18 bl_18 br_18 wl_87 vdd gnd cell_6t
Xbit_r88_c18 bl_18 br_18 wl_88 vdd gnd cell_6t
Xbit_r89_c18 bl_18 br_18 wl_89 vdd gnd cell_6t
Xbit_r90_c18 bl_18 br_18 wl_90 vdd gnd cell_6t
Xbit_r91_c18 bl_18 br_18 wl_91 vdd gnd cell_6t
Xbit_r92_c18 bl_18 br_18 wl_92 vdd gnd cell_6t
Xbit_r93_c18 bl_18 br_18 wl_93 vdd gnd cell_6t
Xbit_r94_c18 bl_18 br_18 wl_94 vdd gnd cell_6t
Xbit_r95_c18 bl_18 br_18 wl_95 vdd gnd cell_6t
Xbit_r96_c18 bl_18 br_18 wl_96 vdd gnd cell_6t
Xbit_r97_c18 bl_18 br_18 wl_97 vdd gnd cell_6t
Xbit_r98_c18 bl_18 br_18 wl_98 vdd gnd cell_6t
Xbit_r99_c18 bl_18 br_18 wl_99 vdd gnd cell_6t
Xbit_r100_c18 bl_18 br_18 wl_100 vdd gnd cell_6t
Xbit_r101_c18 bl_18 br_18 wl_101 vdd gnd cell_6t
Xbit_r102_c18 bl_18 br_18 wl_102 vdd gnd cell_6t
Xbit_r103_c18 bl_18 br_18 wl_103 vdd gnd cell_6t
Xbit_r104_c18 bl_18 br_18 wl_104 vdd gnd cell_6t
Xbit_r105_c18 bl_18 br_18 wl_105 vdd gnd cell_6t
Xbit_r106_c18 bl_18 br_18 wl_106 vdd gnd cell_6t
Xbit_r107_c18 bl_18 br_18 wl_107 vdd gnd cell_6t
Xbit_r108_c18 bl_18 br_18 wl_108 vdd gnd cell_6t
Xbit_r109_c18 bl_18 br_18 wl_109 vdd gnd cell_6t
Xbit_r110_c18 bl_18 br_18 wl_110 vdd gnd cell_6t
Xbit_r111_c18 bl_18 br_18 wl_111 vdd gnd cell_6t
Xbit_r112_c18 bl_18 br_18 wl_112 vdd gnd cell_6t
Xbit_r113_c18 bl_18 br_18 wl_113 vdd gnd cell_6t
Xbit_r114_c18 bl_18 br_18 wl_114 vdd gnd cell_6t
Xbit_r115_c18 bl_18 br_18 wl_115 vdd gnd cell_6t
Xbit_r116_c18 bl_18 br_18 wl_116 vdd gnd cell_6t
Xbit_r117_c18 bl_18 br_18 wl_117 vdd gnd cell_6t
Xbit_r118_c18 bl_18 br_18 wl_118 vdd gnd cell_6t
Xbit_r119_c18 bl_18 br_18 wl_119 vdd gnd cell_6t
Xbit_r120_c18 bl_18 br_18 wl_120 vdd gnd cell_6t
Xbit_r121_c18 bl_18 br_18 wl_121 vdd gnd cell_6t
Xbit_r122_c18 bl_18 br_18 wl_122 vdd gnd cell_6t
Xbit_r123_c18 bl_18 br_18 wl_123 vdd gnd cell_6t
Xbit_r124_c18 bl_18 br_18 wl_124 vdd gnd cell_6t
Xbit_r125_c18 bl_18 br_18 wl_125 vdd gnd cell_6t
Xbit_r126_c18 bl_18 br_18 wl_126 vdd gnd cell_6t
Xbit_r127_c18 bl_18 br_18 wl_127 vdd gnd cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd cell_6t
Xbit_r1_c19 bl_19 br_19 wl_1 vdd gnd cell_6t
Xbit_r2_c19 bl_19 br_19 wl_2 vdd gnd cell_6t
Xbit_r3_c19 bl_19 br_19 wl_3 vdd gnd cell_6t
Xbit_r4_c19 bl_19 br_19 wl_4 vdd gnd cell_6t
Xbit_r5_c19 bl_19 br_19 wl_5 vdd gnd cell_6t
Xbit_r6_c19 bl_19 br_19 wl_6 vdd gnd cell_6t
Xbit_r7_c19 bl_19 br_19 wl_7 vdd gnd cell_6t
Xbit_r8_c19 bl_19 br_19 wl_8 vdd gnd cell_6t
Xbit_r9_c19 bl_19 br_19 wl_9 vdd gnd cell_6t
Xbit_r10_c19 bl_19 br_19 wl_10 vdd gnd cell_6t
Xbit_r11_c19 bl_19 br_19 wl_11 vdd gnd cell_6t
Xbit_r12_c19 bl_19 br_19 wl_12 vdd gnd cell_6t
Xbit_r13_c19 bl_19 br_19 wl_13 vdd gnd cell_6t
Xbit_r14_c19 bl_19 br_19 wl_14 vdd gnd cell_6t
Xbit_r15_c19 bl_19 br_19 wl_15 vdd gnd cell_6t
Xbit_r16_c19 bl_19 br_19 wl_16 vdd gnd cell_6t
Xbit_r17_c19 bl_19 br_19 wl_17 vdd gnd cell_6t
Xbit_r18_c19 bl_19 br_19 wl_18 vdd gnd cell_6t
Xbit_r19_c19 bl_19 br_19 wl_19 vdd gnd cell_6t
Xbit_r20_c19 bl_19 br_19 wl_20 vdd gnd cell_6t
Xbit_r21_c19 bl_19 br_19 wl_21 vdd gnd cell_6t
Xbit_r22_c19 bl_19 br_19 wl_22 vdd gnd cell_6t
Xbit_r23_c19 bl_19 br_19 wl_23 vdd gnd cell_6t
Xbit_r24_c19 bl_19 br_19 wl_24 vdd gnd cell_6t
Xbit_r25_c19 bl_19 br_19 wl_25 vdd gnd cell_6t
Xbit_r26_c19 bl_19 br_19 wl_26 vdd gnd cell_6t
Xbit_r27_c19 bl_19 br_19 wl_27 vdd gnd cell_6t
Xbit_r28_c19 bl_19 br_19 wl_28 vdd gnd cell_6t
Xbit_r29_c19 bl_19 br_19 wl_29 vdd gnd cell_6t
Xbit_r30_c19 bl_19 br_19 wl_30 vdd gnd cell_6t
Xbit_r31_c19 bl_19 br_19 wl_31 vdd gnd cell_6t
Xbit_r32_c19 bl_19 br_19 wl_32 vdd gnd cell_6t
Xbit_r33_c19 bl_19 br_19 wl_33 vdd gnd cell_6t
Xbit_r34_c19 bl_19 br_19 wl_34 vdd gnd cell_6t
Xbit_r35_c19 bl_19 br_19 wl_35 vdd gnd cell_6t
Xbit_r36_c19 bl_19 br_19 wl_36 vdd gnd cell_6t
Xbit_r37_c19 bl_19 br_19 wl_37 vdd gnd cell_6t
Xbit_r38_c19 bl_19 br_19 wl_38 vdd gnd cell_6t
Xbit_r39_c19 bl_19 br_19 wl_39 vdd gnd cell_6t
Xbit_r40_c19 bl_19 br_19 wl_40 vdd gnd cell_6t
Xbit_r41_c19 bl_19 br_19 wl_41 vdd gnd cell_6t
Xbit_r42_c19 bl_19 br_19 wl_42 vdd gnd cell_6t
Xbit_r43_c19 bl_19 br_19 wl_43 vdd gnd cell_6t
Xbit_r44_c19 bl_19 br_19 wl_44 vdd gnd cell_6t
Xbit_r45_c19 bl_19 br_19 wl_45 vdd gnd cell_6t
Xbit_r46_c19 bl_19 br_19 wl_46 vdd gnd cell_6t
Xbit_r47_c19 bl_19 br_19 wl_47 vdd gnd cell_6t
Xbit_r48_c19 bl_19 br_19 wl_48 vdd gnd cell_6t
Xbit_r49_c19 bl_19 br_19 wl_49 vdd gnd cell_6t
Xbit_r50_c19 bl_19 br_19 wl_50 vdd gnd cell_6t
Xbit_r51_c19 bl_19 br_19 wl_51 vdd gnd cell_6t
Xbit_r52_c19 bl_19 br_19 wl_52 vdd gnd cell_6t
Xbit_r53_c19 bl_19 br_19 wl_53 vdd gnd cell_6t
Xbit_r54_c19 bl_19 br_19 wl_54 vdd gnd cell_6t
Xbit_r55_c19 bl_19 br_19 wl_55 vdd gnd cell_6t
Xbit_r56_c19 bl_19 br_19 wl_56 vdd gnd cell_6t
Xbit_r57_c19 bl_19 br_19 wl_57 vdd gnd cell_6t
Xbit_r58_c19 bl_19 br_19 wl_58 vdd gnd cell_6t
Xbit_r59_c19 bl_19 br_19 wl_59 vdd gnd cell_6t
Xbit_r60_c19 bl_19 br_19 wl_60 vdd gnd cell_6t
Xbit_r61_c19 bl_19 br_19 wl_61 vdd gnd cell_6t
Xbit_r62_c19 bl_19 br_19 wl_62 vdd gnd cell_6t
Xbit_r63_c19 bl_19 br_19 wl_63 vdd gnd cell_6t
Xbit_r64_c19 bl_19 br_19 wl_64 vdd gnd cell_6t
Xbit_r65_c19 bl_19 br_19 wl_65 vdd gnd cell_6t
Xbit_r66_c19 bl_19 br_19 wl_66 vdd gnd cell_6t
Xbit_r67_c19 bl_19 br_19 wl_67 vdd gnd cell_6t
Xbit_r68_c19 bl_19 br_19 wl_68 vdd gnd cell_6t
Xbit_r69_c19 bl_19 br_19 wl_69 vdd gnd cell_6t
Xbit_r70_c19 bl_19 br_19 wl_70 vdd gnd cell_6t
Xbit_r71_c19 bl_19 br_19 wl_71 vdd gnd cell_6t
Xbit_r72_c19 bl_19 br_19 wl_72 vdd gnd cell_6t
Xbit_r73_c19 bl_19 br_19 wl_73 vdd gnd cell_6t
Xbit_r74_c19 bl_19 br_19 wl_74 vdd gnd cell_6t
Xbit_r75_c19 bl_19 br_19 wl_75 vdd gnd cell_6t
Xbit_r76_c19 bl_19 br_19 wl_76 vdd gnd cell_6t
Xbit_r77_c19 bl_19 br_19 wl_77 vdd gnd cell_6t
Xbit_r78_c19 bl_19 br_19 wl_78 vdd gnd cell_6t
Xbit_r79_c19 bl_19 br_19 wl_79 vdd gnd cell_6t
Xbit_r80_c19 bl_19 br_19 wl_80 vdd gnd cell_6t
Xbit_r81_c19 bl_19 br_19 wl_81 vdd gnd cell_6t
Xbit_r82_c19 bl_19 br_19 wl_82 vdd gnd cell_6t
Xbit_r83_c19 bl_19 br_19 wl_83 vdd gnd cell_6t
Xbit_r84_c19 bl_19 br_19 wl_84 vdd gnd cell_6t
Xbit_r85_c19 bl_19 br_19 wl_85 vdd gnd cell_6t
Xbit_r86_c19 bl_19 br_19 wl_86 vdd gnd cell_6t
Xbit_r87_c19 bl_19 br_19 wl_87 vdd gnd cell_6t
Xbit_r88_c19 bl_19 br_19 wl_88 vdd gnd cell_6t
Xbit_r89_c19 bl_19 br_19 wl_89 vdd gnd cell_6t
Xbit_r90_c19 bl_19 br_19 wl_90 vdd gnd cell_6t
Xbit_r91_c19 bl_19 br_19 wl_91 vdd gnd cell_6t
Xbit_r92_c19 bl_19 br_19 wl_92 vdd gnd cell_6t
Xbit_r93_c19 bl_19 br_19 wl_93 vdd gnd cell_6t
Xbit_r94_c19 bl_19 br_19 wl_94 vdd gnd cell_6t
Xbit_r95_c19 bl_19 br_19 wl_95 vdd gnd cell_6t
Xbit_r96_c19 bl_19 br_19 wl_96 vdd gnd cell_6t
Xbit_r97_c19 bl_19 br_19 wl_97 vdd gnd cell_6t
Xbit_r98_c19 bl_19 br_19 wl_98 vdd gnd cell_6t
Xbit_r99_c19 bl_19 br_19 wl_99 vdd gnd cell_6t
Xbit_r100_c19 bl_19 br_19 wl_100 vdd gnd cell_6t
Xbit_r101_c19 bl_19 br_19 wl_101 vdd gnd cell_6t
Xbit_r102_c19 bl_19 br_19 wl_102 vdd gnd cell_6t
Xbit_r103_c19 bl_19 br_19 wl_103 vdd gnd cell_6t
Xbit_r104_c19 bl_19 br_19 wl_104 vdd gnd cell_6t
Xbit_r105_c19 bl_19 br_19 wl_105 vdd gnd cell_6t
Xbit_r106_c19 bl_19 br_19 wl_106 vdd gnd cell_6t
Xbit_r107_c19 bl_19 br_19 wl_107 vdd gnd cell_6t
Xbit_r108_c19 bl_19 br_19 wl_108 vdd gnd cell_6t
Xbit_r109_c19 bl_19 br_19 wl_109 vdd gnd cell_6t
Xbit_r110_c19 bl_19 br_19 wl_110 vdd gnd cell_6t
Xbit_r111_c19 bl_19 br_19 wl_111 vdd gnd cell_6t
Xbit_r112_c19 bl_19 br_19 wl_112 vdd gnd cell_6t
Xbit_r113_c19 bl_19 br_19 wl_113 vdd gnd cell_6t
Xbit_r114_c19 bl_19 br_19 wl_114 vdd gnd cell_6t
Xbit_r115_c19 bl_19 br_19 wl_115 vdd gnd cell_6t
Xbit_r116_c19 bl_19 br_19 wl_116 vdd gnd cell_6t
Xbit_r117_c19 bl_19 br_19 wl_117 vdd gnd cell_6t
Xbit_r118_c19 bl_19 br_19 wl_118 vdd gnd cell_6t
Xbit_r119_c19 bl_19 br_19 wl_119 vdd gnd cell_6t
Xbit_r120_c19 bl_19 br_19 wl_120 vdd gnd cell_6t
Xbit_r121_c19 bl_19 br_19 wl_121 vdd gnd cell_6t
Xbit_r122_c19 bl_19 br_19 wl_122 vdd gnd cell_6t
Xbit_r123_c19 bl_19 br_19 wl_123 vdd gnd cell_6t
Xbit_r124_c19 bl_19 br_19 wl_124 vdd gnd cell_6t
Xbit_r125_c19 bl_19 br_19 wl_125 vdd gnd cell_6t
Xbit_r126_c19 bl_19 br_19 wl_126 vdd gnd cell_6t
Xbit_r127_c19 bl_19 br_19 wl_127 vdd gnd cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd cell_6t
Xbit_r1_c20 bl_20 br_20 wl_1 vdd gnd cell_6t
Xbit_r2_c20 bl_20 br_20 wl_2 vdd gnd cell_6t
Xbit_r3_c20 bl_20 br_20 wl_3 vdd gnd cell_6t
Xbit_r4_c20 bl_20 br_20 wl_4 vdd gnd cell_6t
Xbit_r5_c20 bl_20 br_20 wl_5 vdd gnd cell_6t
Xbit_r6_c20 bl_20 br_20 wl_6 vdd gnd cell_6t
Xbit_r7_c20 bl_20 br_20 wl_7 vdd gnd cell_6t
Xbit_r8_c20 bl_20 br_20 wl_8 vdd gnd cell_6t
Xbit_r9_c20 bl_20 br_20 wl_9 vdd gnd cell_6t
Xbit_r10_c20 bl_20 br_20 wl_10 vdd gnd cell_6t
Xbit_r11_c20 bl_20 br_20 wl_11 vdd gnd cell_6t
Xbit_r12_c20 bl_20 br_20 wl_12 vdd gnd cell_6t
Xbit_r13_c20 bl_20 br_20 wl_13 vdd gnd cell_6t
Xbit_r14_c20 bl_20 br_20 wl_14 vdd gnd cell_6t
Xbit_r15_c20 bl_20 br_20 wl_15 vdd gnd cell_6t
Xbit_r16_c20 bl_20 br_20 wl_16 vdd gnd cell_6t
Xbit_r17_c20 bl_20 br_20 wl_17 vdd gnd cell_6t
Xbit_r18_c20 bl_20 br_20 wl_18 vdd gnd cell_6t
Xbit_r19_c20 bl_20 br_20 wl_19 vdd gnd cell_6t
Xbit_r20_c20 bl_20 br_20 wl_20 vdd gnd cell_6t
Xbit_r21_c20 bl_20 br_20 wl_21 vdd gnd cell_6t
Xbit_r22_c20 bl_20 br_20 wl_22 vdd gnd cell_6t
Xbit_r23_c20 bl_20 br_20 wl_23 vdd gnd cell_6t
Xbit_r24_c20 bl_20 br_20 wl_24 vdd gnd cell_6t
Xbit_r25_c20 bl_20 br_20 wl_25 vdd gnd cell_6t
Xbit_r26_c20 bl_20 br_20 wl_26 vdd gnd cell_6t
Xbit_r27_c20 bl_20 br_20 wl_27 vdd gnd cell_6t
Xbit_r28_c20 bl_20 br_20 wl_28 vdd gnd cell_6t
Xbit_r29_c20 bl_20 br_20 wl_29 vdd gnd cell_6t
Xbit_r30_c20 bl_20 br_20 wl_30 vdd gnd cell_6t
Xbit_r31_c20 bl_20 br_20 wl_31 vdd gnd cell_6t
Xbit_r32_c20 bl_20 br_20 wl_32 vdd gnd cell_6t
Xbit_r33_c20 bl_20 br_20 wl_33 vdd gnd cell_6t
Xbit_r34_c20 bl_20 br_20 wl_34 vdd gnd cell_6t
Xbit_r35_c20 bl_20 br_20 wl_35 vdd gnd cell_6t
Xbit_r36_c20 bl_20 br_20 wl_36 vdd gnd cell_6t
Xbit_r37_c20 bl_20 br_20 wl_37 vdd gnd cell_6t
Xbit_r38_c20 bl_20 br_20 wl_38 vdd gnd cell_6t
Xbit_r39_c20 bl_20 br_20 wl_39 vdd gnd cell_6t
Xbit_r40_c20 bl_20 br_20 wl_40 vdd gnd cell_6t
Xbit_r41_c20 bl_20 br_20 wl_41 vdd gnd cell_6t
Xbit_r42_c20 bl_20 br_20 wl_42 vdd gnd cell_6t
Xbit_r43_c20 bl_20 br_20 wl_43 vdd gnd cell_6t
Xbit_r44_c20 bl_20 br_20 wl_44 vdd gnd cell_6t
Xbit_r45_c20 bl_20 br_20 wl_45 vdd gnd cell_6t
Xbit_r46_c20 bl_20 br_20 wl_46 vdd gnd cell_6t
Xbit_r47_c20 bl_20 br_20 wl_47 vdd gnd cell_6t
Xbit_r48_c20 bl_20 br_20 wl_48 vdd gnd cell_6t
Xbit_r49_c20 bl_20 br_20 wl_49 vdd gnd cell_6t
Xbit_r50_c20 bl_20 br_20 wl_50 vdd gnd cell_6t
Xbit_r51_c20 bl_20 br_20 wl_51 vdd gnd cell_6t
Xbit_r52_c20 bl_20 br_20 wl_52 vdd gnd cell_6t
Xbit_r53_c20 bl_20 br_20 wl_53 vdd gnd cell_6t
Xbit_r54_c20 bl_20 br_20 wl_54 vdd gnd cell_6t
Xbit_r55_c20 bl_20 br_20 wl_55 vdd gnd cell_6t
Xbit_r56_c20 bl_20 br_20 wl_56 vdd gnd cell_6t
Xbit_r57_c20 bl_20 br_20 wl_57 vdd gnd cell_6t
Xbit_r58_c20 bl_20 br_20 wl_58 vdd gnd cell_6t
Xbit_r59_c20 bl_20 br_20 wl_59 vdd gnd cell_6t
Xbit_r60_c20 bl_20 br_20 wl_60 vdd gnd cell_6t
Xbit_r61_c20 bl_20 br_20 wl_61 vdd gnd cell_6t
Xbit_r62_c20 bl_20 br_20 wl_62 vdd gnd cell_6t
Xbit_r63_c20 bl_20 br_20 wl_63 vdd gnd cell_6t
Xbit_r64_c20 bl_20 br_20 wl_64 vdd gnd cell_6t
Xbit_r65_c20 bl_20 br_20 wl_65 vdd gnd cell_6t
Xbit_r66_c20 bl_20 br_20 wl_66 vdd gnd cell_6t
Xbit_r67_c20 bl_20 br_20 wl_67 vdd gnd cell_6t
Xbit_r68_c20 bl_20 br_20 wl_68 vdd gnd cell_6t
Xbit_r69_c20 bl_20 br_20 wl_69 vdd gnd cell_6t
Xbit_r70_c20 bl_20 br_20 wl_70 vdd gnd cell_6t
Xbit_r71_c20 bl_20 br_20 wl_71 vdd gnd cell_6t
Xbit_r72_c20 bl_20 br_20 wl_72 vdd gnd cell_6t
Xbit_r73_c20 bl_20 br_20 wl_73 vdd gnd cell_6t
Xbit_r74_c20 bl_20 br_20 wl_74 vdd gnd cell_6t
Xbit_r75_c20 bl_20 br_20 wl_75 vdd gnd cell_6t
Xbit_r76_c20 bl_20 br_20 wl_76 vdd gnd cell_6t
Xbit_r77_c20 bl_20 br_20 wl_77 vdd gnd cell_6t
Xbit_r78_c20 bl_20 br_20 wl_78 vdd gnd cell_6t
Xbit_r79_c20 bl_20 br_20 wl_79 vdd gnd cell_6t
Xbit_r80_c20 bl_20 br_20 wl_80 vdd gnd cell_6t
Xbit_r81_c20 bl_20 br_20 wl_81 vdd gnd cell_6t
Xbit_r82_c20 bl_20 br_20 wl_82 vdd gnd cell_6t
Xbit_r83_c20 bl_20 br_20 wl_83 vdd gnd cell_6t
Xbit_r84_c20 bl_20 br_20 wl_84 vdd gnd cell_6t
Xbit_r85_c20 bl_20 br_20 wl_85 vdd gnd cell_6t
Xbit_r86_c20 bl_20 br_20 wl_86 vdd gnd cell_6t
Xbit_r87_c20 bl_20 br_20 wl_87 vdd gnd cell_6t
Xbit_r88_c20 bl_20 br_20 wl_88 vdd gnd cell_6t
Xbit_r89_c20 bl_20 br_20 wl_89 vdd gnd cell_6t
Xbit_r90_c20 bl_20 br_20 wl_90 vdd gnd cell_6t
Xbit_r91_c20 bl_20 br_20 wl_91 vdd gnd cell_6t
Xbit_r92_c20 bl_20 br_20 wl_92 vdd gnd cell_6t
Xbit_r93_c20 bl_20 br_20 wl_93 vdd gnd cell_6t
Xbit_r94_c20 bl_20 br_20 wl_94 vdd gnd cell_6t
Xbit_r95_c20 bl_20 br_20 wl_95 vdd gnd cell_6t
Xbit_r96_c20 bl_20 br_20 wl_96 vdd gnd cell_6t
Xbit_r97_c20 bl_20 br_20 wl_97 vdd gnd cell_6t
Xbit_r98_c20 bl_20 br_20 wl_98 vdd gnd cell_6t
Xbit_r99_c20 bl_20 br_20 wl_99 vdd gnd cell_6t
Xbit_r100_c20 bl_20 br_20 wl_100 vdd gnd cell_6t
Xbit_r101_c20 bl_20 br_20 wl_101 vdd gnd cell_6t
Xbit_r102_c20 bl_20 br_20 wl_102 vdd gnd cell_6t
Xbit_r103_c20 bl_20 br_20 wl_103 vdd gnd cell_6t
Xbit_r104_c20 bl_20 br_20 wl_104 vdd gnd cell_6t
Xbit_r105_c20 bl_20 br_20 wl_105 vdd gnd cell_6t
Xbit_r106_c20 bl_20 br_20 wl_106 vdd gnd cell_6t
Xbit_r107_c20 bl_20 br_20 wl_107 vdd gnd cell_6t
Xbit_r108_c20 bl_20 br_20 wl_108 vdd gnd cell_6t
Xbit_r109_c20 bl_20 br_20 wl_109 vdd gnd cell_6t
Xbit_r110_c20 bl_20 br_20 wl_110 vdd gnd cell_6t
Xbit_r111_c20 bl_20 br_20 wl_111 vdd gnd cell_6t
Xbit_r112_c20 bl_20 br_20 wl_112 vdd gnd cell_6t
Xbit_r113_c20 bl_20 br_20 wl_113 vdd gnd cell_6t
Xbit_r114_c20 bl_20 br_20 wl_114 vdd gnd cell_6t
Xbit_r115_c20 bl_20 br_20 wl_115 vdd gnd cell_6t
Xbit_r116_c20 bl_20 br_20 wl_116 vdd gnd cell_6t
Xbit_r117_c20 bl_20 br_20 wl_117 vdd gnd cell_6t
Xbit_r118_c20 bl_20 br_20 wl_118 vdd gnd cell_6t
Xbit_r119_c20 bl_20 br_20 wl_119 vdd gnd cell_6t
Xbit_r120_c20 bl_20 br_20 wl_120 vdd gnd cell_6t
Xbit_r121_c20 bl_20 br_20 wl_121 vdd gnd cell_6t
Xbit_r122_c20 bl_20 br_20 wl_122 vdd gnd cell_6t
Xbit_r123_c20 bl_20 br_20 wl_123 vdd gnd cell_6t
Xbit_r124_c20 bl_20 br_20 wl_124 vdd gnd cell_6t
Xbit_r125_c20 bl_20 br_20 wl_125 vdd gnd cell_6t
Xbit_r126_c20 bl_20 br_20 wl_126 vdd gnd cell_6t
Xbit_r127_c20 bl_20 br_20 wl_127 vdd gnd cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd cell_6t
Xbit_r1_c21 bl_21 br_21 wl_1 vdd gnd cell_6t
Xbit_r2_c21 bl_21 br_21 wl_2 vdd gnd cell_6t
Xbit_r3_c21 bl_21 br_21 wl_3 vdd gnd cell_6t
Xbit_r4_c21 bl_21 br_21 wl_4 vdd gnd cell_6t
Xbit_r5_c21 bl_21 br_21 wl_5 vdd gnd cell_6t
Xbit_r6_c21 bl_21 br_21 wl_6 vdd gnd cell_6t
Xbit_r7_c21 bl_21 br_21 wl_7 vdd gnd cell_6t
Xbit_r8_c21 bl_21 br_21 wl_8 vdd gnd cell_6t
Xbit_r9_c21 bl_21 br_21 wl_9 vdd gnd cell_6t
Xbit_r10_c21 bl_21 br_21 wl_10 vdd gnd cell_6t
Xbit_r11_c21 bl_21 br_21 wl_11 vdd gnd cell_6t
Xbit_r12_c21 bl_21 br_21 wl_12 vdd gnd cell_6t
Xbit_r13_c21 bl_21 br_21 wl_13 vdd gnd cell_6t
Xbit_r14_c21 bl_21 br_21 wl_14 vdd gnd cell_6t
Xbit_r15_c21 bl_21 br_21 wl_15 vdd gnd cell_6t
Xbit_r16_c21 bl_21 br_21 wl_16 vdd gnd cell_6t
Xbit_r17_c21 bl_21 br_21 wl_17 vdd gnd cell_6t
Xbit_r18_c21 bl_21 br_21 wl_18 vdd gnd cell_6t
Xbit_r19_c21 bl_21 br_21 wl_19 vdd gnd cell_6t
Xbit_r20_c21 bl_21 br_21 wl_20 vdd gnd cell_6t
Xbit_r21_c21 bl_21 br_21 wl_21 vdd gnd cell_6t
Xbit_r22_c21 bl_21 br_21 wl_22 vdd gnd cell_6t
Xbit_r23_c21 bl_21 br_21 wl_23 vdd gnd cell_6t
Xbit_r24_c21 bl_21 br_21 wl_24 vdd gnd cell_6t
Xbit_r25_c21 bl_21 br_21 wl_25 vdd gnd cell_6t
Xbit_r26_c21 bl_21 br_21 wl_26 vdd gnd cell_6t
Xbit_r27_c21 bl_21 br_21 wl_27 vdd gnd cell_6t
Xbit_r28_c21 bl_21 br_21 wl_28 vdd gnd cell_6t
Xbit_r29_c21 bl_21 br_21 wl_29 vdd gnd cell_6t
Xbit_r30_c21 bl_21 br_21 wl_30 vdd gnd cell_6t
Xbit_r31_c21 bl_21 br_21 wl_31 vdd gnd cell_6t
Xbit_r32_c21 bl_21 br_21 wl_32 vdd gnd cell_6t
Xbit_r33_c21 bl_21 br_21 wl_33 vdd gnd cell_6t
Xbit_r34_c21 bl_21 br_21 wl_34 vdd gnd cell_6t
Xbit_r35_c21 bl_21 br_21 wl_35 vdd gnd cell_6t
Xbit_r36_c21 bl_21 br_21 wl_36 vdd gnd cell_6t
Xbit_r37_c21 bl_21 br_21 wl_37 vdd gnd cell_6t
Xbit_r38_c21 bl_21 br_21 wl_38 vdd gnd cell_6t
Xbit_r39_c21 bl_21 br_21 wl_39 vdd gnd cell_6t
Xbit_r40_c21 bl_21 br_21 wl_40 vdd gnd cell_6t
Xbit_r41_c21 bl_21 br_21 wl_41 vdd gnd cell_6t
Xbit_r42_c21 bl_21 br_21 wl_42 vdd gnd cell_6t
Xbit_r43_c21 bl_21 br_21 wl_43 vdd gnd cell_6t
Xbit_r44_c21 bl_21 br_21 wl_44 vdd gnd cell_6t
Xbit_r45_c21 bl_21 br_21 wl_45 vdd gnd cell_6t
Xbit_r46_c21 bl_21 br_21 wl_46 vdd gnd cell_6t
Xbit_r47_c21 bl_21 br_21 wl_47 vdd gnd cell_6t
Xbit_r48_c21 bl_21 br_21 wl_48 vdd gnd cell_6t
Xbit_r49_c21 bl_21 br_21 wl_49 vdd gnd cell_6t
Xbit_r50_c21 bl_21 br_21 wl_50 vdd gnd cell_6t
Xbit_r51_c21 bl_21 br_21 wl_51 vdd gnd cell_6t
Xbit_r52_c21 bl_21 br_21 wl_52 vdd gnd cell_6t
Xbit_r53_c21 bl_21 br_21 wl_53 vdd gnd cell_6t
Xbit_r54_c21 bl_21 br_21 wl_54 vdd gnd cell_6t
Xbit_r55_c21 bl_21 br_21 wl_55 vdd gnd cell_6t
Xbit_r56_c21 bl_21 br_21 wl_56 vdd gnd cell_6t
Xbit_r57_c21 bl_21 br_21 wl_57 vdd gnd cell_6t
Xbit_r58_c21 bl_21 br_21 wl_58 vdd gnd cell_6t
Xbit_r59_c21 bl_21 br_21 wl_59 vdd gnd cell_6t
Xbit_r60_c21 bl_21 br_21 wl_60 vdd gnd cell_6t
Xbit_r61_c21 bl_21 br_21 wl_61 vdd gnd cell_6t
Xbit_r62_c21 bl_21 br_21 wl_62 vdd gnd cell_6t
Xbit_r63_c21 bl_21 br_21 wl_63 vdd gnd cell_6t
Xbit_r64_c21 bl_21 br_21 wl_64 vdd gnd cell_6t
Xbit_r65_c21 bl_21 br_21 wl_65 vdd gnd cell_6t
Xbit_r66_c21 bl_21 br_21 wl_66 vdd gnd cell_6t
Xbit_r67_c21 bl_21 br_21 wl_67 vdd gnd cell_6t
Xbit_r68_c21 bl_21 br_21 wl_68 vdd gnd cell_6t
Xbit_r69_c21 bl_21 br_21 wl_69 vdd gnd cell_6t
Xbit_r70_c21 bl_21 br_21 wl_70 vdd gnd cell_6t
Xbit_r71_c21 bl_21 br_21 wl_71 vdd gnd cell_6t
Xbit_r72_c21 bl_21 br_21 wl_72 vdd gnd cell_6t
Xbit_r73_c21 bl_21 br_21 wl_73 vdd gnd cell_6t
Xbit_r74_c21 bl_21 br_21 wl_74 vdd gnd cell_6t
Xbit_r75_c21 bl_21 br_21 wl_75 vdd gnd cell_6t
Xbit_r76_c21 bl_21 br_21 wl_76 vdd gnd cell_6t
Xbit_r77_c21 bl_21 br_21 wl_77 vdd gnd cell_6t
Xbit_r78_c21 bl_21 br_21 wl_78 vdd gnd cell_6t
Xbit_r79_c21 bl_21 br_21 wl_79 vdd gnd cell_6t
Xbit_r80_c21 bl_21 br_21 wl_80 vdd gnd cell_6t
Xbit_r81_c21 bl_21 br_21 wl_81 vdd gnd cell_6t
Xbit_r82_c21 bl_21 br_21 wl_82 vdd gnd cell_6t
Xbit_r83_c21 bl_21 br_21 wl_83 vdd gnd cell_6t
Xbit_r84_c21 bl_21 br_21 wl_84 vdd gnd cell_6t
Xbit_r85_c21 bl_21 br_21 wl_85 vdd gnd cell_6t
Xbit_r86_c21 bl_21 br_21 wl_86 vdd gnd cell_6t
Xbit_r87_c21 bl_21 br_21 wl_87 vdd gnd cell_6t
Xbit_r88_c21 bl_21 br_21 wl_88 vdd gnd cell_6t
Xbit_r89_c21 bl_21 br_21 wl_89 vdd gnd cell_6t
Xbit_r90_c21 bl_21 br_21 wl_90 vdd gnd cell_6t
Xbit_r91_c21 bl_21 br_21 wl_91 vdd gnd cell_6t
Xbit_r92_c21 bl_21 br_21 wl_92 vdd gnd cell_6t
Xbit_r93_c21 bl_21 br_21 wl_93 vdd gnd cell_6t
Xbit_r94_c21 bl_21 br_21 wl_94 vdd gnd cell_6t
Xbit_r95_c21 bl_21 br_21 wl_95 vdd gnd cell_6t
Xbit_r96_c21 bl_21 br_21 wl_96 vdd gnd cell_6t
Xbit_r97_c21 bl_21 br_21 wl_97 vdd gnd cell_6t
Xbit_r98_c21 bl_21 br_21 wl_98 vdd gnd cell_6t
Xbit_r99_c21 bl_21 br_21 wl_99 vdd gnd cell_6t
Xbit_r100_c21 bl_21 br_21 wl_100 vdd gnd cell_6t
Xbit_r101_c21 bl_21 br_21 wl_101 vdd gnd cell_6t
Xbit_r102_c21 bl_21 br_21 wl_102 vdd gnd cell_6t
Xbit_r103_c21 bl_21 br_21 wl_103 vdd gnd cell_6t
Xbit_r104_c21 bl_21 br_21 wl_104 vdd gnd cell_6t
Xbit_r105_c21 bl_21 br_21 wl_105 vdd gnd cell_6t
Xbit_r106_c21 bl_21 br_21 wl_106 vdd gnd cell_6t
Xbit_r107_c21 bl_21 br_21 wl_107 vdd gnd cell_6t
Xbit_r108_c21 bl_21 br_21 wl_108 vdd gnd cell_6t
Xbit_r109_c21 bl_21 br_21 wl_109 vdd gnd cell_6t
Xbit_r110_c21 bl_21 br_21 wl_110 vdd gnd cell_6t
Xbit_r111_c21 bl_21 br_21 wl_111 vdd gnd cell_6t
Xbit_r112_c21 bl_21 br_21 wl_112 vdd gnd cell_6t
Xbit_r113_c21 bl_21 br_21 wl_113 vdd gnd cell_6t
Xbit_r114_c21 bl_21 br_21 wl_114 vdd gnd cell_6t
Xbit_r115_c21 bl_21 br_21 wl_115 vdd gnd cell_6t
Xbit_r116_c21 bl_21 br_21 wl_116 vdd gnd cell_6t
Xbit_r117_c21 bl_21 br_21 wl_117 vdd gnd cell_6t
Xbit_r118_c21 bl_21 br_21 wl_118 vdd gnd cell_6t
Xbit_r119_c21 bl_21 br_21 wl_119 vdd gnd cell_6t
Xbit_r120_c21 bl_21 br_21 wl_120 vdd gnd cell_6t
Xbit_r121_c21 bl_21 br_21 wl_121 vdd gnd cell_6t
Xbit_r122_c21 bl_21 br_21 wl_122 vdd gnd cell_6t
Xbit_r123_c21 bl_21 br_21 wl_123 vdd gnd cell_6t
Xbit_r124_c21 bl_21 br_21 wl_124 vdd gnd cell_6t
Xbit_r125_c21 bl_21 br_21 wl_125 vdd gnd cell_6t
Xbit_r126_c21 bl_21 br_21 wl_126 vdd gnd cell_6t
Xbit_r127_c21 bl_21 br_21 wl_127 vdd gnd cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd cell_6t
Xbit_r1_c22 bl_22 br_22 wl_1 vdd gnd cell_6t
Xbit_r2_c22 bl_22 br_22 wl_2 vdd gnd cell_6t
Xbit_r3_c22 bl_22 br_22 wl_3 vdd gnd cell_6t
Xbit_r4_c22 bl_22 br_22 wl_4 vdd gnd cell_6t
Xbit_r5_c22 bl_22 br_22 wl_5 vdd gnd cell_6t
Xbit_r6_c22 bl_22 br_22 wl_6 vdd gnd cell_6t
Xbit_r7_c22 bl_22 br_22 wl_7 vdd gnd cell_6t
Xbit_r8_c22 bl_22 br_22 wl_8 vdd gnd cell_6t
Xbit_r9_c22 bl_22 br_22 wl_9 vdd gnd cell_6t
Xbit_r10_c22 bl_22 br_22 wl_10 vdd gnd cell_6t
Xbit_r11_c22 bl_22 br_22 wl_11 vdd gnd cell_6t
Xbit_r12_c22 bl_22 br_22 wl_12 vdd gnd cell_6t
Xbit_r13_c22 bl_22 br_22 wl_13 vdd gnd cell_6t
Xbit_r14_c22 bl_22 br_22 wl_14 vdd gnd cell_6t
Xbit_r15_c22 bl_22 br_22 wl_15 vdd gnd cell_6t
Xbit_r16_c22 bl_22 br_22 wl_16 vdd gnd cell_6t
Xbit_r17_c22 bl_22 br_22 wl_17 vdd gnd cell_6t
Xbit_r18_c22 bl_22 br_22 wl_18 vdd gnd cell_6t
Xbit_r19_c22 bl_22 br_22 wl_19 vdd gnd cell_6t
Xbit_r20_c22 bl_22 br_22 wl_20 vdd gnd cell_6t
Xbit_r21_c22 bl_22 br_22 wl_21 vdd gnd cell_6t
Xbit_r22_c22 bl_22 br_22 wl_22 vdd gnd cell_6t
Xbit_r23_c22 bl_22 br_22 wl_23 vdd gnd cell_6t
Xbit_r24_c22 bl_22 br_22 wl_24 vdd gnd cell_6t
Xbit_r25_c22 bl_22 br_22 wl_25 vdd gnd cell_6t
Xbit_r26_c22 bl_22 br_22 wl_26 vdd gnd cell_6t
Xbit_r27_c22 bl_22 br_22 wl_27 vdd gnd cell_6t
Xbit_r28_c22 bl_22 br_22 wl_28 vdd gnd cell_6t
Xbit_r29_c22 bl_22 br_22 wl_29 vdd gnd cell_6t
Xbit_r30_c22 bl_22 br_22 wl_30 vdd gnd cell_6t
Xbit_r31_c22 bl_22 br_22 wl_31 vdd gnd cell_6t
Xbit_r32_c22 bl_22 br_22 wl_32 vdd gnd cell_6t
Xbit_r33_c22 bl_22 br_22 wl_33 vdd gnd cell_6t
Xbit_r34_c22 bl_22 br_22 wl_34 vdd gnd cell_6t
Xbit_r35_c22 bl_22 br_22 wl_35 vdd gnd cell_6t
Xbit_r36_c22 bl_22 br_22 wl_36 vdd gnd cell_6t
Xbit_r37_c22 bl_22 br_22 wl_37 vdd gnd cell_6t
Xbit_r38_c22 bl_22 br_22 wl_38 vdd gnd cell_6t
Xbit_r39_c22 bl_22 br_22 wl_39 vdd gnd cell_6t
Xbit_r40_c22 bl_22 br_22 wl_40 vdd gnd cell_6t
Xbit_r41_c22 bl_22 br_22 wl_41 vdd gnd cell_6t
Xbit_r42_c22 bl_22 br_22 wl_42 vdd gnd cell_6t
Xbit_r43_c22 bl_22 br_22 wl_43 vdd gnd cell_6t
Xbit_r44_c22 bl_22 br_22 wl_44 vdd gnd cell_6t
Xbit_r45_c22 bl_22 br_22 wl_45 vdd gnd cell_6t
Xbit_r46_c22 bl_22 br_22 wl_46 vdd gnd cell_6t
Xbit_r47_c22 bl_22 br_22 wl_47 vdd gnd cell_6t
Xbit_r48_c22 bl_22 br_22 wl_48 vdd gnd cell_6t
Xbit_r49_c22 bl_22 br_22 wl_49 vdd gnd cell_6t
Xbit_r50_c22 bl_22 br_22 wl_50 vdd gnd cell_6t
Xbit_r51_c22 bl_22 br_22 wl_51 vdd gnd cell_6t
Xbit_r52_c22 bl_22 br_22 wl_52 vdd gnd cell_6t
Xbit_r53_c22 bl_22 br_22 wl_53 vdd gnd cell_6t
Xbit_r54_c22 bl_22 br_22 wl_54 vdd gnd cell_6t
Xbit_r55_c22 bl_22 br_22 wl_55 vdd gnd cell_6t
Xbit_r56_c22 bl_22 br_22 wl_56 vdd gnd cell_6t
Xbit_r57_c22 bl_22 br_22 wl_57 vdd gnd cell_6t
Xbit_r58_c22 bl_22 br_22 wl_58 vdd gnd cell_6t
Xbit_r59_c22 bl_22 br_22 wl_59 vdd gnd cell_6t
Xbit_r60_c22 bl_22 br_22 wl_60 vdd gnd cell_6t
Xbit_r61_c22 bl_22 br_22 wl_61 vdd gnd cell_6t
Xbit_r62_c22 bl_22 br_22 wl_62 vdd gnd cell_6t
Xbit_r63_c22 bl_22 br_22 wl_63 vdd gnd cell_6t
Xbit_r64_c22 bl_22 br_22 wl_64 vdd gnd cell_6t
Xbit_r65_c22 bl_22 br_22 wl_65 vdd gnd cell_6t
Xbit_r66_c22 bl_22 br_22 wl_66 vdd gnd cell_6t
Xbit_r67_c22 bl_22 br_22 wl_67 vdd gnd cell_6t
Xbit_r68_c22 bl_22 br_22 wl_68 vdd gnd cell_6t
Xbit_r69_c22 bl_22 br_22 wl_69 vdd gnd cell_6t
Xbit_r70_c22 bl_22 br_22 wl_70 vdd gnd cell_6t
Xbit_r71_c22 bl_22 br_22 wl_71 vdd gnd cell_6t
Xbit_r72_c22 bl_22 br_22 wl_72 vdd gnd cell_6t
Xbit_r73_c22 bl_22 br_22 wl_73 vdd gnd cell_6t
Xbit_r74_c22 bl_22 br_22 wl_74 vdd gnd cell_6t
Xbit_r75_c22 bl_22 br_22 wl_75 vdd gnd cell_6t
Xbit_r76_c22 bl_22 br_22 wl_76 vdd gnd cell_6t
Xbit_r77_c22 bl_22 br_22 wl_77 vdd gnd cell_6t
Xbit_r78_c22 bl_22 br_22 wl_78 vdd gnd cell_6t
Xbit_r79_c22 bl_22 br_22 wl_79 vdd gnd cell_6t
Xbit_r80_c22 bl_22 br_22 wl_80 vdd gnd cell_6t
Xbit_r81_c22 bl_22 br_22 wl_81 vdd gnd cell_6t
Xbit_r82_c22 bl_22 br_22 wl_82 vdd gnd cell_6t
Xbit_r83_c22 bl_22 br_22 wl_83 vdd gnd cell_6t
Xbit_r84_c22 bl_22 br_22 wl_84 vdd gnd cell_6t
Xbit_r85_c22 bl_22 br_22 wl_85 vdd gnd cell_6t
Xbit_r86_c22 bl_22 br_22 wl_86 vdd gnd cell_6t
Xbit_r87_c22 bl_22 br_22 wl_87 vdd gnd cell_6t
Xbit_r88_c22 bl_22 br_22 wl_88 vdd gnd cell_6t
Xbit_r89_c22 bl_22 br_22 wl_89 vdd gnd cell_6t
Xbit_r90_c22 bl_22 br_22 wl_90 vdd gnd cell_6t
Xbit_r91_c22 bl_22 br_22 wl_91 vdd gnd cell_6t
Xbit_r92_c22 bl_22 br_22 wl_92 vdd gnd cell_6t
Xbit_r93_c22 bl_22 br_22 wl_93 vdd gnd cell_6t
Xbit_r94_c22 bl_22 br_22 wl_94 vdd gnd cell_6t
Xbit_r95_c22 bl_22 br_22 wl_95 vdd gnd cell_6t
Xbit_r96_c22 bl_22 br_22 wl_96 vdd gnd cell_6t
Xbit_r97_c22 bl_22 br_22 wl_97 vdd gnd cell_6t
Xbit_r98_c22 bl_22 br_22 wl_98 vdd gnd cell_6t
Xbit_r99_c22 bl_22 br_22 wl_99 vdd gnd cell_6t
Xbit_r100_c22 bl_22 br_22 wl_100 vdd gnd cell_6t
Xbit_r101_c22 bl_22 br_22 wl_101 vdd gnd cell_6t
Xbit_r102_c22 bl_22 br_22 wl_102 vdd gnd cell_6t
Xbit_r103_c22 bl_22 br_22 wl_103 vdd gnd cell_6t
Xbit_r104_c22 bl_22 br_22 wl_104 vdd gnd cell_6t
Xbit_r105_c22 bl_22 br_22 wl_105 vdd gnd cell_6t
Xbit_r106_c22 bl_22 br_22 wl_106 vdd gnd cell_6t
Xbit_r107_c22 bl_22 br_22 wl_107 vdd gnd cell_6t
Xbit_r108_c22 bl_22 br_22 wl_108 vdd gnd cell_6t
Xbit_r109_c22 bl_22 br_22 wl_109 vdd gnd cell_6t
Xbit_r110_c22 bl_22 br_22 wl_110 vdd gnd cell_6t
Xbit_r111_c22 bl_22 br_22 wl_111 vdd gnd cell_6t
Xbit_r112_c22 bl_22 br_22 wl_112 vdd gnd cell_6t
Xbit_r113_c22 bl_22 br_22 wl_113 vdd gnd cell_6t
Xbit_r114_c22 bl_22 br_22 wl_114 vdd gnd cell_6t
Xbit_r115_c22 bl_22 br_22 wl_115 vdd gnd cell_6t
Xbit_r116_c22 bl_22 br_22 wl_116 vdd gnd cell_6t
Xbit_r117_c22 bl_22 br_22 wl_117 vdd gnd cell_6t
Xbit_r118_c22 bl_22 br_22 wl_118 vdd gnd cell_6t
Xbit_r119_c22 bl_22 br_22 wl_119 vdd gnd cell_6t
Xbit_r120_c22 bl_22 br_22 wl_120 vdd gnd cell_6t
Xbit_r121_c22 bl_22 br_22 wl_121 vdd gnd cell_6t
Xbit_r122_c22 bl_22 br_22 wl_122 vdd gnd cell_6t
Xbit_r123_c22 bl_22 br_22 wl_123 vdd gnd cell_6t
Xbit_r124_c22 bl_22 br_22 wl_124 vdd gnd cell_6t
Xbit_r125_c22 bl_22 br_22 wl_125 vdd gnd cell_6t
Xbit_r126_c22 bl_22 br_22 wl_126 vdd gnd cell_6t
Xbit_r127_c22 bl_22 br_22 wl_127 vdd gnd cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd cell_6t
Xbit_r1_c23 bl_23 br_23 wl_1 vdd gnd cell_6t
Xbit_r2_c23 bl_23 br_23 wl_2 vdd gnd cell_6t
Xbit_r3_c23 bl_23 br_23 wl_3 vdd gnd cell_6t
Xbit_r4_c23 bl_23 br_23 wl_4 vdd gnd cell_6t
Xbit_r5_c23 bl_23 br_23 wl_5 vdd gnd cell_6t
Xbit_r6_c23 bl_23 br_23 wl_6 vdd gnd cell_6t
Xbit_r7_c23 bl_23 br_23 wl_7 vdd gnd cell_6t
Xbit_r8_c23 bl_23 br_23 wl_8 vdd gnd cell_6t
Xbit_r9_c23 bl_23 br_23 wl_9 vdd gnd cell_6t
Xbit_r10_c23 bl_23 br_23 wl_10 vdd gnd cell_6t
Xbit_r11_c23 bl_23 br_23 wl_11 vdd gnd cell_6t
Xbit_r12_c23 bl_23 br_23 wl_12 vdd gnd cell_6t
Xbit_r13_c23 bl_23 br_23 wl_13 vdd gnd cell_6t
Xbit_r14_c23 bl_23 br_23 wl_14 vdd gnd cell_6t
Xbit_r15_c23 bl_23 br_23 wl_15 vdd gnd cell_6t
Xbit_r16_c23 bl_23 br_23 wl_16 vdd gnd cell_6t
Xbit_r17_c23 bl_23 br_23 wl_17 vdd gnd cell_6t
Xbit_r18_c23 bl_23 br_23 wl_18 vdd gnd cell_6t
Xbit_r19_c23 bl_23 br_23 wl_19 vdd gnd cell_6t
Xbit_r20_c23 bl_23 br_23 wl_20 vdd gnd cell_6t
Xbit_r21_c23 bl_23 br_23 wl_21 vdd gnd cell_6t
Xbit_r22_c23 bl_23 br_23 wl_22 vdd gnd cell_6t
Xbit_r23_c23 bl_23 br_23 wl_23 vdd gnd cell_6t
Xbit_r24_c23 bl_23 br_23 wl_24 vdd gnd cell_6t
Xbit_r25_c23 bl_23 br_23 wl_25 vdd gnd cell_6t
Xbit_r26_c23 bl_23 br_23 wl_26 vdd gnd cell_6t
Xbit_r27_c23 bl_23 br_23 wl_27 vdd gnd cell_6t
Xbit_r28_c23 bl_23 br_23 wl_28 vdd gnd cell_6t
Xbit_r29_c23 bl_23 br_23 wl_29 vdd gnd cell_6t
Xbit_r30_c23 bl_23 br_23 wl_30 vdd gnd cell_6t
Xbit_r31_c23 bl_23 br_23 wl_31 vdd gnd cell_6t
Xbit_r32_c23 bl_23 br_23 wl_32 vdd gnd cell_6t
Xbit_r33_c23 bl_23 br_23 wl_33 vdd gnd cell_6t
Xbit_r34_c23 bl_23 br_23 wl_34 vdd gnd cell_6t
Xbit_r35_c23 bl_23 br_23 wl_35 vdd gnd cell_6t
Xbit_r36_c23 bl_23 br_23 wl_36 vdd gnd cell_6t
Xbit_r37_c23 bl_23 br_23 wl_37 vdd gnd cell_6t
Xbit_r38_c23 bl_23 br_23 wl_38 vdd gnd cell_6t
Xbit_r39_c23 bl_23 br_23 wl_39 vdd gnd cell_6t
Xbit_r40_c23 bl_23 br_23 wl_40 vdd gnd cell_6t
Xbit_r41_c23 bl_23 br_23 wl_41 vdd gnd cell_6t
Xbit_r42_c23 bl_23 br_23 wl_42 vdd gnd cell_6t
Xbit_r43_c23 bl_23 br_23 wl_43 vdd gnd cell_6t
Xbit_r44_c23 bl_23 br_23 wl_44 vdd gnd cell_6t
Xbit_r45_c23 bl_23 br_23 wl_45 vdd gnd cell_6t
Xbit_r46_c23 bl_23 br_23 wl_46 vdd gnd cell_6t
Xbit_r47_c23 bl_23 br_23 wl_47 vdd gnd cell_6t
Xbit_r48_c23 bl_23 br_23 wl_48 vdd gnd cell_6t
Xbit_r49_c23 bl_23 br_23 wl_49 vdd gnd cell_6t
Xbit_r50_c23 bl_23 br_23 wl_50 vdd gnd cell_6t
Xbit_r51_c23 bl_23 br_23 wl_51 vdd gnd cell_6t
Xbit_r52_c23 bl_23 br_23 wl_52 vdd gnd cell_6t
Xbit_r53_c23 bl_23 br_23 wl_53 vdd gnd cell_6t
Xbit_r54_c23 bl_23 br_23 wl_54 vdd gnd cell_6t
Xbit_r55_c23 bl_23 br_23 wl_55 vdd gnd cell_6t
Xbit_r56_c23 bl_23 br_23 wl_56 vdd gnd cell_6t
Xbit_r57_c23 bl_23 br_23 wl_57 vdd gnd cell_6t
Xbit_r58_c23 bl_23 br_23 wl_58 vdd gnd cell_6t
Xbit_r59_c23 bl_23 br_23 wl_59 vdd gnd cell_6t
Xbit_r60_c23 bl_23 br_23 wl_60 vdd gnd cell_6t
Xbit_r61_c23 bl_23 br_23 wl_61 vdd gnd cell_6t
Xbit_r62_c23 bl_23 br_23 wl_62 vdd gnd cell_6t
Xbit_r63_c23 bl_23 br_23 wl_63 vdd gnd cell_6t
Xbit_r64_c23 bl_23 br_23 wl_64 vdd gnd cell_6t
Xbit_r65_c23 bl_23 br_23 wl_65 vdd gnd cell_6t
Xbit_r66_c23 bl_23 br_23 wl_66 vdd gnd cell_6t
Xbit_r67_c23 bl_23 br_23 wl_67 vdd gnd cell_6t
Xbit_r68_c23 bl_23 br_23 wl_68 vdd gnd cell_6t
Xbit_r69_c23 bl_23 br_23 wl_69 vdd gnd cell_6t
Xbit_r70_c23 bl_23 br_23 wl_70 vdd gnd cell_6t
Xbit_r71_c23 bl_23 br_23 wl_71 vdd gnd cell_6t
Xbit_r72_c23 bl_23 br_23 wl_72 vdd gnd cell_6t
Xbit_r73_c23 bl_23 br_23 wl_73 vdd gnd cell_6t
Xbit_r74_c23 bl_23 br_23 wl_74 vdd gnd cell_6t
Xbit_r75_c23 bl_23 br_23 wl_75 vdd gnd cell_6t
Xbit_r76_c23 bl_23 br_23 wl_76 vdd gnd cell_6t
Xbit_r77_c23 bl_23 br_23 wl_77 vdd gnd cell_6t
Xbit_r78_c23 bl_23 br_23 wl_78 vdd gnd cell_6t
Xbit_r79_c23 bl_23 br_23 wl_79 vdd gnd cell_6t
Xbit_r80_c23 bl_23 br_23 wl_80 vdd gnd cell_6t
Xbit_r81_c23 bl_23 br_23 wl_81 vdd gnd cell_6t
Xbit_r82_c23 bl_23 br_23 wl_82 vdd gnd cell_6t
Xbit_r83_c23 bl_23 br_23 wl_83 vdd gnd cell_6t
Xbit_r84_c23 bl_23 br_23 wl_84 vdd gnd cell_6t
Xbit_r85_c23 bl_23 br_23 wl_85 vdd gnd cell_6t
Xbit_r86_c23 bl_23 br_23 wl_86 vdd gnd cell_6t
Xbit_r87_c23 bl_23 br_23 wl_87 vdd gnd cell_6t
Xbit_r88_c23 bl_23 br_23 wl_88 vdd gnd cell_6t
Xbit_r89_c23 bl_23 br_23 wl_89 vdd gnd cell_6t
Xbit_r90_c23 bl_23 br_23 wl_90 vdd gnd cell_6t
Xbit_r91_c23 bl_23 br_23 wl_91 vdd gnd cell_6t
Xbit_r92_c23 bl_23 br_23 wl_92 vdd gnd cell_6t
Xbit_r93_c23 bl_23 br_23 wl_93 vdd gnd cell_6t
Xbit_r94_c23 bl_23 br_23 wl_94 vdd gnd cell_6t
Xbit_r95_c23 bl_23 br_23 wl_95 vdd gnd cell_6t
Xbit_r96_c23 bl_23 br_23 wl_96 vdd gnd cell_6t
Xbit_r97_c23 bl_23 br_23 wl_97 vdd gnd cell_6t
Xbit_r98_c23 bl_23 br_23 wl_98 vdd gnd cell_6t
Xbit_r99_c23 bl_23 br_23 wl_99 vdd gnd cell_6t
Xbit_r100_c23 bl_23 br_23 wl_100 vdd gnd cell_6t
Xbit_r101_c23 bl_23 br_23 wl_101 vdd gnd cell_6t
Xbit_r102_c23 bl_23 br_23 wl_102 vdd gnd cell_6t
Xbit_r103_c23 bl_23 br_23 wl_103 vdd gnd cell_6t
Xbit_r104_c23 bl_23 br_23 wl_104 vdd gnd cell_6t
Xbit_r105_c23 bl_23 br_23 wl_105 vdd gnd cell_6t
Xbit_r106_c23 bl_23 br_23 wl_106 vdd gnd cell_6t
Xbit_r107_c23 bl_23 br_23 wl_107 vdd gnd cell_6t
Xbit_r108_c23 bl_23 br_23 wl_108 vdd gnd cell_6t
Xbit_r109_c23 bl_23 br_23 wl_109 vdd gnd cell_6t
Xbit_r110_c23 bl_23 br_23 wl_110 vdd gnd cell_6t
Xbit_r111_c23 bl_23 br_23 wl_111 vdd gnd cell_6t
Xbit_r112_c23 bl_23 br_23 wl_112 vdd gnd cell_6t
Xbit_r113_c23 bl_23 br_23 wl_113 vdd gnd cell_6t
Xbit_r114_c23 bl_23 br_23 wl_114 vdd gnd cell_6t
Xbit_r115_c23 bl_23 br_23 wl_115 vdd gnd cell_6t
Xbit_r116_c23 bl_23 br_23 wl_116 vdd gnd cell_6t
Xbit_r117_c23 bl_23 br_23 wl_117 vdd gnd cell_6t
Xbit_r118_c23 bl_23 br_23 wl_118 vdd gnd cell_6t
Xbit_r119_c23 bl_23 br_23 wl_119 vdd gnd cell_6t
Xbit_r120_c23 bl_23 br_23 wl_120 vdd gnd cell_6t
Xbit_r121_c23 bl_23 br_23 wl_121 vdd gnd cell_6t
Xbit_r122_c23 bl_23 br_23 wl_122 vdd gnd cell_6t
Xbit_r123_c23 bl_23 br_23 wl_123 vdd gnd cell_6t
Xbit_r124_c23 bl_23 br_23 wl_124 vdd gnd cell_6t
Xbit_r125_c23 bl_23 br_23 wl_125 vdd gnd cell_6t
Xbit_r126_c23 bl_23 br_23 wl_126 vdd gnd cell_6t
Xbit_r127_c23 bl_23 br_23 wl_127 vdd gnd cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd cell_6t
Xbit_r1_c24 bl_24 br_24 wl_1 vdd gnd cell_6t
Xbit_r2_c24 bl_24 br_24 wl_2 vdd gnd cell_6t
Xbit_r3_c24 bl_24 br_24 wl_3 vdd gnd cell_6t
Xbit_r4_c24 bl_24 br_24 wl_4 vdd gnd cell_6t
Xbit_r5_c24 bl_24 br_24 wl_5 vdd gnd cell_6t
Xbit_r6_c24 bl_24 br_24 wl_6 vdd gnd cell_6t
Xbit_r7_c24 bl_24 br_24 wl_7 vdd gnd cell_6t
Xbit_r8_c24 bl_24 br_24 wl_8 vdd gnd cell_6t
Xbit_r9_c24 bl_24 br_24 wl_9 vdd gnd cell_6t
Xbit_r10_c24 bl_24 br_24 wl_10 vdd gnd cell_6t
Xbit_r11_c24 bl_24 br_24 wl_11 vdd gnd cell_6t
Xbit_r12_c24 bl_24 br_24 wl_12 vdd gnd cell_6t
Xbit_r13_c24 bl_24 br_24 wl_13 vdd gnd cell_6t
Xbit_r14_c24 bl_24 br_24 wl_14 vdd gnd cell_6t
Xbit_r15_c24 bl_24 br_24 wl_15 vdd gnd cell_6t
Xbit_r16_c24 bl_24 br_24 wl_16 vdd gnd cell_6t
Xbit_r17_c24 bl_24 br_24 wl_17 vdd gnd cell_6t
Xbit_r18_c24 bl_24 br_24 wl_18 vdd gnd cell_6t
Xbit_r19_c24 bl_24 br_24 wl_19 vdd gnd cell_6t
Xbit_r20_c24 bl_24 br_24 wl_20 vdd gnd cell_6t
Xbit_r21_c24 bl_24 br_24 wl_21 vdd gnd cell_6t
Xbit_r22_c24 bl_24 br_24 wl_22 vdd gnd cell_6t
Xbit_r23_c24 bl_24 br_24 wl_23 vdd gnd cell_6t
Xbit_r24_c24 bl_24 br_24 wl_24 vdd gnd cell_6t
Xbit_r25_c24 bl_24 br_24 wl_25 vdd gnd cell_6t
Xbit_r26_c24 bl_24 br_24 wl_26 vdd gnd cell_6t
Xbit_r27_c24 bl_24 br_24 wl_27 vdd gnd cell_6t
Xbit_r28_c24 bl_24 br_24 wl_28 vdd gnd cell_6t
Xbit_r29_c24 bl_24 br_24 wl_29 vdd gnd cell_6t
Xbit_r30_c24 bl_24 br_24 wl_30 vdd gnd cell_6t
Xbit_r31_c24 bl_24 br_24 wl_31 vdd gnd cell_6t
Xbit_r32_c24 bl_24 br_24 wl_32 vdd gnd cell_6t
Xbit_r33_c24 bl_24 br_24 wl_33 vdd gnd cell_6t
Xbit_r34_c24 bl_24 br_24 wl_34 vdd gnd cell_6t
Xbit_r35_c24 bl_24 br_24 wl_35 vdd gnd cell_6t
Xbit_r36_c24 bl_24 br_24 wl_36 vdd gnd cell_6t
Xbit_r37_c24 bl_24 br_24 wl_37 vdd gnd cell_6t
Xbit_r38_c24 bl_24 br_24 wl_38 vdd gnd cell_6t
Xbit_r39_c24 bl_24 br_24 wl_39 vdd gnd cell_6t
Xbit_r40_c24 bl_24 br_24 wl_40 vdd gnd cell_6t
Xbit_r41_c24 bl_24 br_24 wl_41 vdd gnd cell_6t
Xbit_r42_c24 bl_24 br_24 wl_42 vdd gnd cell_6t
Xbit_r43_c24 bl_24 br_24 wl_43 vdd gnd cell_6t
Xbit_r44_c24 bl_24 br_24 wl_44 vdd gnd cell_6t
Xbit_r45_c24 bl_24 br_24 wl_45 vdd gnd cell_6t
Xbit_r46_c24 bl_24 br_24 wl_46 vdd gnd cell_6t
Xbit_r47_c24 bl_24 br_24 wl_47 vdd gnd cell_6t
Xbit_r48_c24 bl_24 br_24 wl_48 vdd gnd cell_6t
Xbit_r49_c24 bl_24 br_24 wl_49 vdd gnd cell_6t
Xbit_r50_c24 bl_24 br_24 wl_50 vdd gnd cell_6t
Xbit_r51_c24 bl_24 br_24 wl_51 vdd gnd cell_6t
Xbit_r52_c24 bl_24 br_24 wl_52 vdd gnd cell_6t
Xbit_r53_c24 bl_24 br_24 wl_53 vdd gnd cell_6t
Xbit_r54_c24 bl_24 br_24 wl_54 vdd gnd cell_6t
Xbit_r55_c24 bl_24 br_24 wl_55 vdd gnd cell_6t
Xbit_r56_c24 bl_24 br_24 wl_56 vdd gnd cell_6t
Xbit_r57_c24 bl_24 br_24 wl_57 vdd gnd cell_6t
Xbit_r58_c24 bl_24 br_24 wl_58 vdd gnd cell_6t
Xbit_r59_c24 bl_24 br_24 wl_59 vdd gnd cell_6t
Xbit_r60_c24 bl_24 br_24 wl_60 vdd gnd cell_6t
Xbit_r61_c24 bl_24 br_24 wl_61 vdd gnd cell_6t
Xbit_r62_c24 bl_24 br_24 wl_62 vdd gnd cell_6t
Xbit_r63_c24 bl_24 br_24 wl_63 vdd gnd cell_6t
Xbit_r64_c24 bl_24 br_24 wl_64 vdd gnd cell_6t
Xbit_r65_c24 bl_24 br_24 wl_65 vdd gnd cell_6t
Xbit_r66_c24 bl_24 br_24 wl_66 vdd gnd cell_6t
Xbit_r67_c24 bl_24 br_24 wl_67 vdd gnd cell_6t
Xbit_r68_c24 bl_24 br_24 wl_68 vdd gnd cell_6t
Xbit_r69_c24 bl_24 br_24 wl_69 vdd gnd cell_6t
Xbit_r70_c24 bl_24 br_24 wl_70 vdd gnd cell_6t
Xbit_r71_c24 bl_24 br_24 wl_71 vdd gnd cell_6t
Xbit_r72_c24 bl_24 br_24 wl_72 vdd gnd cell_6t
Xbit_r73_c24 bl_24 br_24 wl_73 vdd gnd cell_6t
Xbit_r74_c24 bl_24 br_24 wl_74 vdd gnd cell_6t
Xbit_r75_c24 bl_24 br_24 wl_75 vdd gnd cell_6t
Xbit_r76_c24 bl_24 br_24 wl_76 vdd gnd cell_6t
Xbit_r77_c24 bl_24 br_24 wl_77 vdd gnd cell_6t
Xbit_r78_c24 bl_24 br_24 wl_78 vdd gnd cell_6t
Xbit_r79_c24 bl_24 br_24 wl_79 vdd gnd cell_6t
Xbit_r80_c24 bl_24 br_24 wl_80 vdd gnd cell_6t
Xbit_r81_c24 bl_24 br_24 wl_81 vdd gnd cell_6t
Xbit_r82_c24 bl_24 br_24 wl_82 vdd gnd cell_6t
Xbit_r83_c24 bl_24 br_24 wl_83 vdd gnd cell_6t
Xbit_r84_c24 bl_24 br_24 wl_84 vdd gnd cell_6t
Xbit_r85_c24 bl_24 br_24 wl_85 vdd gnd cell_6t
Xbit_r86_c24 bl_24 br_24 wl_86 vdd gnd cell_6t
Xbit_r87_c24 bl_24 br_24 wl_87 vdd gnd cell_6t
Xbit_r88_c24 bl_24 br_24 wl_88 vdd gnd cell_6t
Xbit_r89_c24 bl_24 br_24 wl_89 vdd gnd cell_6t
Xbit_r90_c24 bl_24 br_24 wl_90 vdd gnd cell_6t
Xbit_r91_c24 bl_24 br_24 wl_91 vdd gnd cell_6t
Xbit_r92_c24 bl_24 br_24 wl_92 vdd gnd cell_6t
Xbit_r93_c24 bl_24 br_24 wl_93 vdd gnd cell_6t
Xbit_r94_c24 bl_24 br_24 wl_94 vdd gnd cell_6t
Xbit_r95_c24 bl_24 br_24 wl_95 vdd gnd cell_6t
Xbit_r96_c24 bl_24 br_24 wl_96 vdd gnd cell_6t
Xbit_r97_c24 bl_24 br_24 wl_97 vdd gnd cell_6t
Xbit_r98_c24 bl_24 br_24 wl_98 vdd gnd cell_6t
Xbit_r99_c24 bl_24 br_24 wl_99 vdd gnd cell_6t
Xbit_r100_c24 bl_24 br_24 wl_100 vdd gnd cell_6t
Xbit_r101_c24 bl_24 br_24 wl_101 vdd gnd cell_6t
Xbit_r102_c24 bl_24 br_24 wl_102 vdd gnd cell_6t
Xbit_r103_c24 bl_24 br_24 wl_103 vdd gnd cell_6t
Xbit_r104_c24 bl_24 br_24 wl_104 vdd gnd cell_6t
Xbit_r105_c24 bl_24 br_24 wl_105 vdd gnd cell_6t
Xbit_r106_c24 bl_24 br_24 wl_106 vdd gnd cell_6t
Xbit_r107_c24 bl_24 br_24 wl_107 vdd gnd cell_6t
Xbit_r108_c24 bl_24 br_24 wl_108 vdd gnd cell_6t
Xbit_r109_c24 bl_24 br_24 wl_109 vdd gnd cell_6t
Xbit_r110_c24 bl_24 br_24 wl_110 vdd gnd cell_6t
Xbit_r111_c24 bl_24 br_24 wl_111 vdd gnd cell_6t
Xbit_r112_c24 bl_24 br_24 wl_112 vdd gnd cell_6t
Xbit_r113_c24 bl_24 br_24 wl_113 vdd gnd cell_6t
Xbit_r114_c24 bl_24 br_24 wl_114 vdd gnd cell_6t
Xbit_r115_c24 bl_24 br_24 wl_115 vdd gnd cell_6t
Xbit_r116_c24 bl_24 br_24 wl_116 vdd gnd cell_6t
Xbit_r117_c24 bl_24 br_24 wl_117 vdd gnd cell_6t
Xbit_r118_c24 bl_24 br_24 wl_118 vdd gnd cell_6t
Xbit_r119_c24 bl_24 br_24 wl_119 vdd gnd cell_6t
Xbit_r120_c24 bl_24 br_24 wl_120 vdd gnd cell_6t
Xbit_r121_c24 bl_24 br_24 wl_121 vdd gnd cell_6t
Xbit_r122_c24 bl_24 br_24 wl_122 vdd gnd cell_6t
Xbit_r123_c24 bl_24 br_24 wl_123 vdd gnd cell_6t
Xbit_r124_c24 bl_24 br_24 wl_124 vdd gnd cell_6t
Xbit_r125_c24 bl_24 br_24 wl_125 vdd gnd cell_6t
Xbit_r126_c24 bl_24 br_24 wl_126 vdd gnd cell_6t
Xbit_r127_c24 bl_24 br_24 wl_127 vdd gnd cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd cell_6t
Xbit_r1_c25 bl_25 br_25 wl_1 vdd gnd cell_6t
Xbit_r2_c25 bl_25 br_25 wl_2 vdd gnd cell_6t
Xbit_r3_c25 bl_25 br_25 wl_3 vdd gnd cell_6t
Xbit_r4_c25 bl_25 br_25 wl_4 vdd gnd cell_6t
Xbit_r5_c25 bl_25 br_25 wl_5 vdd gnd cell_6t
Xbit_r6_c25 bl_25 br_25 wl_6 vdd gnd cell_6t
Xbit_r7_c25 bl_25 br_25 wl_7 vdd gnd cell_6t
Xbit_r8_c25 bl_25 br_25 wl_8 vdd gnd cell_6t
Xbit_r9_c25 bl_25 br_25 wl_9 vdd gnd cell_6t
Xbit_r10_c25 bl_25 br_25 wl_10 vdd gnd cell_6t
Xbit_r11_c25 bl_25 br_25 wl_11 vdd gnd cell_6t
Xbit_r12_c25 bl_25 br_25 wl_12 vdd gnd cell_6t
Xbit_r13_c25 bl_25 br_25 wl_13 vdd gnd cell_6t
Xbit_r14_c25 bl_25 br_25 wl_14 vdd gnd cell_6t
Xbit_r15_c25 bl_25 br_25 wl_15 vdd gnd cell_6t
Xbit_r16_c25 bl_25 br_25 wl_16 vdd gnd cell_6t
Xbit_r17_c25 bl_25 br_25 wl_17 vdd gnd cell_6t
Xbit_r18_c25 bl_25 br_25 wl_18 vdd gnd cell_6t
Xbit_r19_c25 bl_25 br_25 wl_19 vdd gnd cell_6t
Xbit_r20_c25 bl_25 br_25 wl_20 vdd gnd cell_6t
Xbit_r21_c25 bl_25 br_25 wl_21 vdd gnd cell_6t
Xbit_r22_c25 bl_25 br_25 wl_22 vdd gnd cell_6t
Xbit_r23_c25 bl_25 br_25 wl_23 vdd gnd cell_6t
Xbit_r24_c25 bl_25 br_25 wl_24 vdd gnd cell_6t
Xbit_r25_c25 bl_25 br_25 wl_25 vdd gnd cell_6t
Xbit_r26_c25 bl_25 br_25 wl_26 vdd gnd cell_6t
Xbit_r27_c25 bl_25 br_25 wl_27 vdd gnd cell_6t
Xbit_r28_c25 bl_25 br_25 wl_28 vdd gnd cell_6t
Xbit_r29_c25 bl_25 br_25 wl_29 vdd gnd cell_6t
Xbit_r30_c25 bl_25 br_25 wl_30 vdd gnd cell_6t
Xbit_r31_c25 bl_25 br_25 wl_31 vdd gnd cell_6t
Xbit_r32_c25 bl_25 br_25 wl_32 vdd gnd cell_6t
Xbit_r33_c25 bl_25 br_25 wl_33 vdd gnd cell_6t
Xbit_r34_c25 bl_25 br_25 wl_34 vdd gnd cell_6t
Xbit_r35_c25 bl_25 br_25 wl_35 vdd gnd cell_6t
Xbit_r36_c25 bl_25 br_25 wl_36 vdd gnd cell_6t
Xbit_r37_c25 bl_25 br_25 wl_37 vdd gnd cell_6t
Xbit_r38_c25 bl_25 br_25 wl_38 vdd gnd cell_6t
Xbit_r39_c25 bl_25 br_25 wl_39 vdd gnd cell_6t
Xbit_r40_c25 bl_25 br_25 wl_40 vdd gnd cell_6t
Xbit_r41_c25 bl_25 br_25 wl_41 vdd gnd cell_6t
Xbit_r42_c25 bl_25 br_25 wl_42 vdd gnd cell_6t
Xbit_r43_c25 bl_25 br_25 wl_43 vdd gnd cell_6t
Xbit_r44_c25 bl_25 br_25 wl_44 vdd gnd cell_6t
Xbit_r45_c25 bl_25 br_25 wl_45 vdd gnd cell_6t
Xbit_r46_c25 bl_25 br_25 wl_46 vdd gnd cell_6t
Xbit_r47_c25 bl_25 br_25 wl_47 vdd gnd cell_6t
Xbit_r48_c25 bl_25 br_25 wl_48 vdd gnd cell_6t
Xbit_r49_c25 bl_25 br_25 wl_49 vdd gnd cell_6t
Xbit_r50_c25 bl_25 br_25 wl_50 vdd gnd cell_6t
Xbit_r51_c25 bl_25 br_25 wl_51 vdd gnd cell_6t
Xbit_r52_c25 bl_25 br_25 wl_52 vdd gnd cell_6t
Xbit_r53_c25 bl_25 br_25 wl_53 vdd gnd cell_6t
Xbit_r54_c25 bl_25 br_25 wl_54 vdd gnd cell_6t
Xbit_r55_c25 bl_25 br_25 wl_55 vdd gnd cell_6t
Xbit_r56_c25 bl_25 br_25 wl_56 vdd gnd cell_6t
Xbit_r57_c25 bl_25 br_25 wl_57 vdd gnd cell_6t
Xbit_r58_c25 bl_25 br_25 wl_58 vdd gnd cell_6t
Xbit_r59_c25 bl_25 br_25 wl_59 vdd gnd cell_6t
Xbit_r60_c25 bl_25 br_25 wl_60 vdd gnd cell_6t
Xbit_r61_c25 bl_25 br_25 wl_61 vdd gnd cell_6t
Xbit_r62_c25 bl_25 br_25 wl_62 vdd gnd cell_6t
Xbit_r63_c25 bl_25 br_25 wl_63 vdd gnd cell_6t
Xbit_r64_c25 bl_25 br_25 wl_64 vdd gnd cell_6t
Xbit_r65_c25 bl_25 br_25 wl_65 vdd gnd cell_6t
Xbit_r66_c25 bl_25 br_25 wl_66 vdd gnd cell_6t
Xbit_r67_c25 bl_25 br_25 wl_67 vdd gnd cell_6t
Xbit_r68_c25 bl_25 br_25 wl_68 vdd gnd cell_6t
Xbit_r69_c25 bl_25 br_25 wl_69 vdd gnd cell_6t
Xbit_r70_c25 bl_25 br_25 wl_70 vdd gnd cell_6t
Xbit_r71_c25 bl_25 br_25 wl_71 vdd gnd cell_6t
Xbit_r72_c25 bl_25 br_25 wl_72 vdd gnd cell_6t
Xbit_r73_c25 bl_25 br_25 wl_73 vdd gnd cell_6t
Xbit_r74_c25 bl_25 br_25 wl_74 vdd gnd cell_6t
Xbit_r75_c25 bl_25 br_25 wl_75 vdd gnd cell_6t
Xbit_r76_c25 bl_25 br_25 wl_76 vdd gnd cell_6t
Xbit_r77_c25 bl_25 br_25 wl_77 vdd gnd cell_6t
Xbit_r78_c25 bl_25 br_25 wl_78 vdd gnd cell_6t
Xbit_r79_c25 bl_25 br_25 wl_79 vdd gnd cell_6t
Xbit_r80_c25 bl_25 br_25 wl_80 vdd gnd cell_6t
Xbit_r81_c25 bl_25 br_25 wl_81 vdd gnd cell_6t
Xbit_r82_c25 bl_25 br_25 wl_82 vdd gnd cell_6t
Xbit_r83_c25 bl_25 br_25 wl_83 vdd gnd cell_6t
Xbit_r84_c25 bl_25 br_25 wl_84 vdd gnd cell_6t
Xbit_r85_c25 bl_25 br_25 wl_85 vdd gnd cell_6t
Xbit_r86_c25 bl_25 br_25 wl_86 vdd gnd cell_6t
Xbit_r87_c25 bl_25 br_25 wl_87 vdd gnd cell_6t
Xbit_r88_c25 bl_25 br_25 wl_88 vdd gnd cell_6t
Xbit_r89_c25 bl_25 br_25 wl_89 vdd gnd cell_6t
Xbit_r90_c25 bl_25 br_25 wl_90 vdd gnd cell_6t
Xbit_r91_c25 bl_25 br_25 wl_91 vdd gnd cell_6t
Xbit_r92_c25 bl_25 br_25 wl_92 vdd gnd cell_6t
Xbit_r93_c25 bl_25 br_25 wl_93 vdd gnd cell_6t
Xbit_r94_c25 bl_25 br_25 wl_94 vdd gnd cell_6t
Xbit_r95_c25 bl_25 br_25 wl_95 vdd gnd cell_6t
Xbit_r96_c25 bl_25 br_25 wl_96 vdd gnd cell_6t
Xbit_r97_c25 bl_25 br_25 wl_97 vdd gnd cell_6t
Xbit_r98_c25 bl_25 br_25 wl_98 vdd gnd cell_6t
Xbit_r99_c25 bl_25 br_25 wl_99 vdd gnd cell_6t
Xbit_r100_c25 bl_25 br_25 wl_100 vdd gnd cell_6t
Xbit_r101_c25 bl_25 br_25 wl_101 vdd gnd cell_6t
Xbit_r102_c25 bl_25 br_25 wl_102 vdd gnd cell_6t
Xbit_r103_c25 bl_25 br_25 wl_103 vdd gnd cell_6t
Xbit_r104_c25 bl_25 br_25 wl_104 vdd gnd cell_6t
Xbit_r105_c25 bl_25 br_25 wl_105 vdd gnd cell_6t
Xbit_r106_c25 bl_25 br_25 wl_106 vdd gnd cell_6t
Xbit_r107_c25 bl_25 br_25 wl_107 vdd gnd cell_6t
Xbit_r108_c25 bl_25 br_25 wl_108 vdd gnd cell_6t
Xbit_r109_c25 bl_25 br_25 wl_109 vdd gnd cell_6t
Xbit_r110_c25 bl_25 br_25 wl_110 vdd gnd cell_6t
Xbit_r111_c25 bl_25 br_25 wl_111 vdd gnd cell_6t
Xbit_r112_c25 bl_25 br_25 wl_112 vdd gnd cell_6t
Xbit_r113_c25 bl_25 br_25 wl_113 vdd gnd cell_6t
Xbit_r114_c25 bl_25 br_25 wl_114 vdd gnd cell_6t
Xbit_r115_c25 bl_25 br_25 wl_115 vdd gnd cell_6t
Xbit_r116_c25 bl_25 br_25 wl_116 vdd gnd cell_6t
Xbit_r117_c25 bl_25 br_25 wl_117 vdd gnd cell_6t
Xbit_r118_c25 bl_25 br_25 wl_118 vdd gnd cell_6t
Xbit_r119_c25 bl_25 br_25 wl_119 vdd gnd cell_6t
Xbit_r120_c25 bl_25 br_25 wl_120 vdd gnd cell_6t
Xbit_r121_c25 bl_25 br_25 wl_121 vdd gnd cell_6t
Xbit_r122_c25 bl_25 br_25 wl_122 vdd gnd cell_6t
Xbit_r123_c25 bl_25 br_25 wl_123 vdd gnd cell_6t
Xbit_r124_c25 bl_25 br_25 wl_124 vdd gnd cell_6t
Xbit_r125_c25 bl_25 br_25 wl_125 vdd gnd cell_6t
Xbit_r126_c25 bl_25 br_25 wl_126 vdd gnd cell_6t
Xbit_r127_c25 bl_25 br_25 wl_127 vdd gnd cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd cell_6t
Xbit_r1_c26 bl_26 br_26 wl_1 vdd gnd cell_6t
Xbit_r2_c26 bl_26 br_26 wl_2 vdd gnd cell_6t
Xbit_r3_c26 bl_26 br_26 wl_3 vdd gnd cell_6t
Xbit_r4_c26 bl_26 br_26 wl_4 vdd gnd cell_6t
Xbit_r5_c26 bl_26 br_26 wl_5 vdd gnd cell_6t
Xbit_r6_c26 bl_26 br_26 wl_6 vdd gnd cell_6t
Xbit_r7_c26 bl_26 br_26 wl_7 vdd gnd cell_6t
Xbit_r8_c26 bl_26 br_26 wl_8 vdd gnd cell_6t
Xbit_r9_c26 bl_26 br_26 wl_9 vdd gnd cell_6t
Xbit_r10_c26 bl_26 br_26 wl_10 vdd gnd cell_6t
Xbit_r11_c26 bl_26 br_26 wl_11 vdd gnd cell_6t
Xbit_r12_c26 bl_26 br_26 wl_12 vdd gnd cell_6t
Xbit_r13_c26 bl_26 br_26 wl_13 vdd gnd cell_6t
Xbit_r14_c26 bl_26 br_26 wl_14 vdd gnd cell_6t
Xbit_r15_c26 bl_26 br_26 wl_15 vdd gnd cell_6t
Xbit_r16_c26 bl_26 br_26 wl_16 vdd gnd cell_6t
Xbit_r17_c26 bl_26 br_26 wl_17 vdd gnd cell_6t
Xbit_r18_c26 bl_26 br_26 wl_18 vdd gnd cell_6t
Xbit_r19_c26 bl_26 br_26 wl_19 vdd gnd cell_6t
Xbit_r20_c26 bl_26 br_26 wl_20 vdd gnd cell_6t
Xbit_r21_c26 bl_26 br_26 wl_21 vdd gnd cell_6t
Xbit_r22_c26 bl_26 br_26 wl_22 vdd gnd cell_6t
Xbit_r23_c26 bl_26 br_26 wl_23 vdd gnd cell_6t
Xbit_r24_c26 bl_26 br_26 wl_24 vdd gnd cell_6t
Xbit_r25_c26 bl_26 br_26 wl_25 vdd gnd cell_6t
Xbit_r26_c26 bl_26 br_26 wl_26 vdd gnd cell_6t
Xbit_r27_c26 bl_26 br_26 wl_27 vdd gnd cell_6t
Xbit_r28_c26 bl_26 br_26 wl_28 vdd gnd cell_6t
Xbit_r29_c26 bl_26 br_26 wl_29 vdd gnd cell_6t
Xbit_r30_c26 bl_26 br_26 wl_30 vdd gnd cell_6t
Xbit_r31_c26 bl_26 br_26 wl_31 vdd gnd cell_6t
Xbit_r32_c26 bl_26 br_26 wl_32 vdd gnd cell_6t
Xbit_r33_c26 bl_26 br_26 wl_33 vdd gnd cell_6t
Xbit_r34_c26 bl_26 br_26 wl_34 vdd gnd cell_6t
Xbit_r35_c26 bl_26 br_26 wl_35 vdd gnd cell_6t
Xbit_r36_c26 bl_26 br_26 wl_36 vdd gnd cell_6t
Xbit_r37_c26 bl_26 br_26 wl_37 vdd gnd cell_6t
Xbit_r38_c26 bl_26 br_26 wl_38 vdd gnd cell_6t
Xbit_r39_c26 bl_26 br_26 wl_39 vdd gnd cell_6t
Xbit_r40_c26 bl_26 br_26 wl_40 vdd gnd cell_6t
Xbit_r41_c26 bl_26 br_26 wl_41 vdd gnd cell_6t
Xbit_r42_c26 bl_26 br_26 wl_42 vdd gnd cell_6t
Xbit_r43_c26 bl_26 br_26 wl_43 vdd gnd cell_6t
Xbit_r44_c26 bl_26 br_26 wl_44 vdd gnd cell_6t
Xbit_r45_c26 bl_26 br_26 wl_45 vdd gnd cell_6t
Xbit_r46_c26 bl_26 br_26 wl_46 vdd gnd cell_6t
Xbit_r47_c26 bl_26 br_26 wl_47 vdd gnd cell_6t
Xbit_r48_c26 bl_26 br_26 wl_48 vdd gnd cell_6t
Xbit_r49_c26 bl_26 br_26 wl_49 vdd gnd cell_6t
Xbit_r50_c26 bl_26 br_26 wl_50 vdd gnd cell_6t
Xbit_r51_c26 bl_26 br_26 wl_51 vdd gnd cell_6t
Xbit_r52_c26 bl_26 br_26 wl_52 vdd gnd cell_6t
Xbit_r53_c26 bl_26 br_26 wl_53 vdd gnd cell_6t
Xbit_r54_c26 bl_26 br_26 wl_54 vdd gnd cell_6t
Xbit_r55_c26 bl_26 br_26 wl_55 vdd gnd cell_6t
Xbit_r56_c26 bl_26 br_26 wl_56 vdd gnd cell_6t
Xbit_r57_c26 bl_26 br_26 wl_57 vdd gnd cell_6t
Xbit_r58_c26 bl_26 br_26 wl_58 vdd gnd cell_6t
Xbit_r59_c26 bl_26 br_26 wl_59 vdd gnd cell_6t
Xbit_r60_c26 bl_26 br_26 wl_60 vdd gnd cell_6t
Xbit_r61_c26 bl_26 br_26 wl_61 vdd gnd cell_6t
Xbit_r62_c26 bl_26 br_26 wl_62 vdd gnd cell_6t
Xbit_r63_c26 bl_26 br_26 wl_63 vdd gnd cell_6t
Xbit_r64_c26 bl_26 br_26 wl_64 vdd gnd cell_6t
Xbit_r65_c26 bl_26 br_26 wl_65 vdd gnd cell_6t
Xbit_r66_c26 bl_26 br_26 wl_66 vdd gnd cell_6t
Xbit_r67_c26 bl_26 br_26 wl_67 vdd gnd cell_6t
Xbit_r68_c26 bl_26 br_26 wl_68 vdd gnd cell_6t
Xbit_r69_c26 bl_26 br_26 wl_69 vdd gnd cell_6t
Xbit_r70_c26 bl_26 br_26 wl_70 vdd gnd cell_6t
Xbit_r71_c26 bl_26 br_26 wl_71 vdd gnd cell_6t
Xbit_r72_c26 bl_26 br_26 wl_72 vdd gnd cell_6t
Xbit_r73_c26 bl_26 br_26 wl_73 vdd gnd cell_6t
Xbit_r74_c26 bl_26 br_26 wl_74 vdd gnd cell_6t
Xbit_r75_c26 bl_26 br_26 wl_75 vdd gnd cell_6t
Xbit_r76_c26 bl_26 br_26 wl_76 vdd gnd cell_6t
Xbit_r77_c26 bl_26 br_26 wl_77 vdd gnd cell_6t
Xbit_r78_c26 bl_26 br_26 wl_78 vdd gnd cell_6t
Xbit_r79_c26 bl_26 br_26 wl_79 vdd gnd cell_6t
Xbit_r80_c26 bl_26 br_26 wl_80 vdd gnd cell_6t
Xbit_r81_c26 bl_26 br_26 wl_81 vdd gnd cell_6t
Xbit_r82_c26 bl_26 br_26 wl_82 vdd gnd cell_6t
Xbit_r83_c26 bl_26 br_26 wl_83 vdd gnd cell_6t
Xbit_r84_c26 bl_26 br_26 wl_84 vdd gnd cell_6t
Xbit_r85_c26 bl_26 br_26 wl_85 vdd gnd cell_6t
Xbit_r86_c26 bl_26 br_26 wl_86 vdd gnd cell_6t
Xbit_r87_c26 bl_26 br_26 wl_87 vdd gnd cell_6t
Xbit_r88_c26 bl_26 br_26 wl_88 vdd gnd cell_6t
Xbit_r89_c26 bl_26 br_26 wl_89 vdd gnd cell_6t
Xbit_r90_c26 bl_26 br_26 wl_90 vdd gnd cell_6t
Xbit_r91_c26 bl_26 br_26 wl_91 vdd gnd cell_6t
Xbit_r92_c26 bl_26 br_26 wl_92 vdd gnd cell_6t
Xbit_r93_c26 bl_26 br_26 wl_93 vdd gnd cell_6t
Xbit_r94_c26 bl_26 br_26 wl_94 vdd gnd cell_6t
Xbit_r95_c26 bl_26 br_26 wl_95 vdd gnd cell_6t
Xbit_r96_c26 bl_26 br_26 wl_96 vdd gnd cell_6t
Xbit_r97_c26 bl_26 br_26 wl_97 vdd gnd cell_6t
Xbit_r98_c26 bl_26 br_26 wl_98 vdd gnd cell_6t
Xbit_r99_c26 bl_26 br_26 wl_99 vdd gnd cell_6t
Xbit_r100_c26 bl_26 br_26 wl_100 vdd gnd cell_6t
Xbit_r101_c26 bl_26 br_26 wl_101 vdd gnd cell_6t
Xbit_r102_c26 bl_26 br_26 wl_102 vdd gnd cell_6t
Xbit_r103_c26 bl_26 br_26 wl_103 vdd gnd cell_6t
Xbit_r104_c26 bl_26 br_26 wl_104 vdd gnd cell_6t
Xbit_r105_c26 bl_26 br_26 wl_105 vdd gnd cell_6t
Xbit_r106_c26 bl_26 br_26 wl_106 vdd gnd cell_6t
Xbit_r107_c26 bl_26 br_26 wl_107 vdd gnd cell_6t
Xbit_r108_c26 bl_26 br_26 wl_108 vdd gnd cell_6t
Xbit_r109_c26 bl_26 br_26 wl_109 vdd gnd cell_6t
Xbit_r110_c26 bl_26 br_26 wl_110 vdd gnd cell_6t
Xbit_r111_c26 bl_26 br_26 wl_111 vdd gnd cell_6t
Xbit_r112_c26 bl_26 br_26 wl_112 vdd gnd cell_6t
Xbit_r113_c26 bl_26 br_26 wl_113 vdd gnd cell_6t
Xbit_r114_c26 bl_26 br_26 wl_114 vdd gnd cell_6t
Xbit_r115_c26 bl_26 br_26 wl_115 vdd gnd cell_6t
Xbit_r116_c26 bl_26 br_26 wl_116 vdd gnd cell_6t
Xbit_r117_c26 bl_26 br_26 wl_117 vdd gnd cell_6t
Xbit_r118_c26 bl_26 br_26 wl_118 vdd gnd cell_6t
Xbit_r119_c26 bl_26 br_26 wl_119 vdd gnd cell_6t
Xbit_r120_c26 bl_26 br_26 wl_120 vdd gnd cell_6t
Xbit_r121_c26 bl_26 br_26 wl_121 vdd gnd cell_6t
Xbit_r122_c26 bl_26 br_26 wl_122 vdd gnd cell_6t
Xbit_r123_c26 bl_26 br_26 wl_123 vdd gnd cell_6t
Xbit_r124_c26 bl_26 br_26 wl_124 vdd gnd cell_6t
Xbit_r125_c26 bl_26 br_26 wl_125 vdd gnd cell_6t
Xbit_r126_c26 bl_26 br_26 wl_126 vdd gnd cell_6t
Xbit_r127_c26 bl_26 br_26 wl_127 vdd gnd cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd cell_6t
Xbit_r1_c27 bl_27 br_27 wl_1 vdd gnd cell_6t
Xbit_r2_c27 bl_27 br_27 wl_2 vdd gnd cell_6t
Xbit_r3_c27 bl_27 br_27 wl_3 vdd gnd cell_6t
Xbit_r4_c27 bl_27 br_27 wl_4 vdd gnd cell_6t
Xbit_r5_c27 bl_27 br_27 wl_5 vdd gnd cell_6t
Xbit_r6_c27 bl_27 br_27 wl_6 vdd gnd cell_6t
Xbit_r7_c27 bl_27 br_27 wl_7 vdd gnd cell_6t
Xbit_r8_c27 bl_27 br_27 wl_8 vdd gnd cell_6t
Xbit_r9_c27 bl_27 br_27 wl_9 vdd gnd cell_6t
Xbit_r10_c27 bl_27 br_27 wl_10 vdd gnd cell_6t
Xbit_r11_c27 bl_27 br_27 wl_11 vdd gnd cell_6t
Xbit_r12_c27 bl_27 br_27 wl_12 vdd gnd cell_6t
Xbit_r13_c27 bl_27 br_27 wl_13 vdd gnd cell_6t
Xbit_r14_c27 bl_27 br_27 wl_14 vdd gnd cell_6t
Xbit_r15_c27 bl_27 br_27 wl_15 vdd gnd cell_6t
Xbit_r16_c27 bl_27 br_27 wl_16 vdd gnd cell_6t
Xbit_r17_c27 bl_27 br_27 wl_17 vdd gnd cell_6t
Xbit_r18_c27 bl_27 br_27 wl_18 vdd gnd cell_6t
Xbit_r19_c27 bl_27 br_27 wl_19 vdd gnd cell_6t
Xbit_r20_c27 bl_27 br_27 wl_20 vdd gnd cell_6t
Xbit_r21_c27 bl_27 br_27 wl_21 vdd gnd cell_6t
Xbit_r22_c27 bl_27 br_27 wl_22 vdd gnd cell_6t
Xbit_r23_c27 bl_27 br_27 wl_23 vdd gnd cell_6t
Xbit_r24_c27 bl_27 br_27 wl_24 vdd gnd cell_6t
Xbit_r25_c27 bl_27 br_27 wl_25 vdd gnd cell_6t
Xbit_r26_c27 bl_27 br_27 wl_26 vdd gnd cell_6t
Xbit_r27_c27 bl_27 br_27 wl_27 vdd gnd cell_6t
Xbit_r28_c27 bl_27 br_27 wl_28 vdd gnd cell_6t
Xbit_r29_c27 bl_27 br_27 wl_29 vdd gnd cell_6t
Xbit_r30_c27 bl_27 br_27 wl_30 vdd gnd cell_6t
Xbit_r31_c27 bl_27 br_27 wl_31 vdd gnd cell_6t
Xbit_r32_c27 bl_27 br_27 wl_32 vdd gnd cell_6t
Xbit_r33_c27 bl_27 br_27 wl_33 vdd gnd cell_6t
Xbit_r34_c27 bl_27 br_27 wl_34 vdd gnd cell_6t
Xbit_r35_c27 bl_27 br_27 wl_35 vdd gnd cell_6t
Xbit_r36_c27 bl_27 br_27 wl_36 vdd gnd cell_6t
Xbit_r37_c27 bl_27 br_27 wl_37 vdd gnd cell_6t
Xbit_r38_c27 bl_27 br_27 wl_38 vdd gnd cell_6t
Xbit_r39_c27 bl_27 br_27 wl_39 vdd gnd cell_6t
Xbit_r40_c27 bl_27 br_27 wl_40 vdd gnd cell_6t
Xbit_r41_c27 bl_27 br_27 wl_41 vdd gnd cell_6t
Xbit_r42_c27 bl_27 br_27 wl_42 vdd gnd cell_6t
Xbit_r43_c27 bl_27 br_27 wl_43 vdd gnd cell_6t
Xbit_r44_c27 bl_27 br_27 wl_44 vdd gnd cell_6t
Xbit_r45_c27 bl_27 br_27 wl_45 vdd gnd cell_6t
Xbit_r46_c27 bl_27 br_27 wl_46 vdd gnd cell_6t
Xbit_r47_c27 bl_27 br_27 wl_47 vdd gnd cell_6t
Xbit_r48_c27 bl_27 br_27 wl_48 vdd gnd cell_6t
Xbit_r49_c27 bl_27 br_27 wl_49 vdd gnd cell_6t
Xbit_r50_c27 bl_27 br_27 wl_50 vdd gnd cell_6t
Xbit_r51_c27 bl_27 br_27 wl_51 vdd gnd cell_6t
Xbit_r52_c27 bl_27 br_27 wl_52 vdd gnd cell_6t
Xbit_r53_c27 bl_27 br_27 wl_53 vdd gnd cell_6t
Xbit_r54_c27 bl_27 br_27 wl_54 vdd gnd cell_6t
Xbit_r55_c27 bl_27 br_27 wl_55 vdd gnd cell_6t
Xbit_r56_c27 bl_27 br_27 wl_56 vdd gnd cell_6t
Xbit_r57_c27 bl_27 br_27 wl_57 vdd gnd cell_6t
Xbit_r58_c27 bl_27 br_27 wl_58 vdd gnd cell_6t
Xbit_r59_c27 bl_27 br_27 wl_59 vdd gnd cell_6t
Xbit_r60_c27 bl_27 br_27 wl_60 vdd gnd cell_6t
Xbit_r61_c27 bl_27 br_27 wl_61 vdd gnd cell_6t
Xbit_r62_c27 bl_27 br_27 wl_62 vdd gnd cell_6t
Xbit_r63_c27 bl_27 br_27 wl_63 vdd gnd cell_6t
Xbit_r64_c27 bl_27 br_27 wl_64 vdd gnd cell_6t
Xbit_r65_c27 bl_27 br_27 wl_65 vdd gnd cell_6t
Xbit_r66_c27 bl_27 br_27 wl_66 vdd gnd cell_6t
Xbit_r67_c27 bl_27 br_27 wl_67 vdd gnd cell_6t
Xbit_r68_c27 bl_27 br_27 wl_68 vdd gnd cell_6t
Xbit_r69_c27 bl_27 br_27 wl_69 vdd gnd cell_6t
Xbit_r70_c27 bl_27 br_27 wl_70 vdd gnd cell_6t
Xbit_r71_c27 bl_27 br_27 wl_71 vdd gnd cell_6t
Xbit_r72_c27 bl_27 br_27 wl_72 vdd gnd cell_6t
Xbit_r73_c27 bl_27 br_27 wl_73 vdd gnd cell_6t
Xbit_r74_c27 bl_27 br_27 wl_74 vdd gnd cell_6t
Xbit_r75_c27 bl_27 br_27 wl_75 vdd gnd cell_6t
Xbit_r76_c27 bl_27 br_27 wl_76 vdd gnd cell_6t
Xbit_r77_c27 bl_27 br_27 wl_77 vdd gnd cell_6t
Xbit_r78_c27 bl_27 br_27 wl_78 vdd gnd cell_6t
Xbit_r79_c27 bl_27 br_27 wl_79 vdd gnd cell_6t
Xbit_r80_c27 bl_27 br_27 wl_80 vdd gnd cell_6t
Xbit_r81_c27 bl_27 br_27 wl_81 vdd gnd cell_6t
Xbit_r82_c27 bl_27 br_27 wl_82 vdd gnd cell_6t
Xbit_r83_c27 bl_27 br_27 wl_83 vdd gnd cell_6t
Xbit_r84_c27 bl_27 br_27 wl_84 vdd gnd cell_6t
Xbit_r85_c27 bl_27 br_27 wl_85 vdd gnd cell_6t
Xbit_r86_c27 bl_27 br_27 wl_86 vdd gnd cell_6t
Xbit_r87_c27 bl_27 br_27 wl_87 vdd gnd cell_6t
Xbit_r88_c27 bl_27 br_27 wl_88 vdd gnd cell_6t
Xbit_r89_c27 bl_27 br_27 wl_89 vdd gnd cell_6t
Xbit_r90_c27 bl_27 br_27 wl_90 vdd gnd cell_6t
Xbit_r91_c27 bl_27 br_27 wl_91 vdd gnd cell_6t
Xbit_r92_c27 bl_27 br_27 wl_92 vdd gnd cell_6t
Xbit_r93_c27 bl_27 br_27 wl_93 vdd gnd cell_6t
Xbit_r94_c27 bl_27 br_27 wl_94 vdd gnd cell_6t
Xbit_r95_c27 bl_27 br_27 wl_95 vdd gnd cell_6t
Xbit_r96_c27 bl_27 br_27 wl_96 vdd gnd cell_6t
Xbit_r97_c27 bl_27 br_27 wl_97 vdd gnd cell_6t
Xbit_r98_c27 bl_27 br_27 wl_98 vdd gnd cell_6t
Xbit_r99_c27 bl_27 br_27 wl_99 vdd gnd cell_6t
Xbit_r100_c27 bl_27 br_27 wl_100 vdd gnd cell_6t
Xbit_r101_c27 bl_27 br_27 wl_101 vdd gnd cell_6t
Xbit_r102_c27 bl_27 br_27 wl_102 vdd gnd cell_6t
Xbit_r103_c27 bl_27 br_27 wl_103 vdd gnd cell_6t
Xbit_r104_c27 bl_27 br_27 wl_104 vdd gnd cell_6t
Xbit_r105_c27 bl_27 br_27 wl_105 vdd gnd cell_6t
Xbit_r106_c27 bl_27 br_27 wl_106 vdd gnd cell_6t
Xbit_r107_c27 bl_27 br_27 wl_107 vdd gnd cell_6t
Xbit_r108_c27 bl_27 br_27 wl_108 vdd gnd cell_6t
Xbit_r109_c27 bl_27 br_27 wl_109 vdd gnd cell_6t
Xbit_r110_c27 bl_27 br_27 wl_110 vdd gnd cell_6t
Xbit_r111_c27 bl_27 br_27 wl_111 vdd gnd cell_6t
Xbit_r112_c27 bl_27 br_27 wl_112 vdd gnd cell_6t
Xbit_r113_c27 bl_27 br_27 wl_113 vdd gnd cell_6t
Xbit_r114_c27 bl_27 br_27 wl_114 vdd gnd cell_6t
Xbit_r115_c27 bl_27 br_27 wl_115 vdd gnd cell_6t
Xbit_r116_c27 bl_27 br_27 wl_116 vdd gnd cell_6t
Xbit_r117_c27 bl_27 br_27 wl_117 vdd gnd cell_6t
Xbit_r118_c27 bl_27 br_27 wl_118 vdd gnd cell_6t
Xbit_r119_c27 bl_27 br_27 wl_119 vdd gnd cell_6t
Xbit_r120_c27 bl_27 br_27 wl_120 vdd gnd cell_6t
Xbit_r121_c27 bl_27 br_27 wl_121 vdd gnd cell_6t
Xbit_r122_c27 bl_27 br_27 wl_122 vdd gnd cell_6t
Xbit_r123_c27 bl_27 br_27 wl_123 vdd gnd cell_6t
Xbit_r124_c27 bl_27 br_27 wl_124 vdd gnd cell_6t
Xbit_r125_c27 bl_27 br_27 wl_125 vdd gnd cell_6t
Xbit_r126_c27 bl_27 br_27 wl_126 vdd gnd cell_6t
Xbit_r127_c27 bl_27 br_27 wl_127 vdd gnd cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd cell_6t
Xbit_r1_c28 bl_28 br_28 wl_1 vdd gnd cell_6t
Xbit_r2_c28 bl_28 br_28 wl_2 vdd gnd cell_6t
Xbit_r3_c28 bl_28 br_28 wl_3 vdd gnd cell_6t
Xbit_r4_c28 bl_28 br_28 wl_4 vdd gnd cell_6t
Xbit_r5_c28 bl_28 br_28 wl_5 vdd gnd cell_6t
Xbit_r6_c28 bl_28 br_28 wl_6 vdd gnd cell_6t
Xbit_r7_c28 bl_28 br_28 wl_7 vdd gnd cell_6t
Xbit_r8_c28 bl_28 br_28 wl_8 vdd gnd cell_6t
Xbit_r9_c28 bl_28 br_28 wl_9 vdd gnd cell_6t
Xbit_r10_c28 bl_28 br_28 wl_10 vdd gnd cell_6t
Xbit_r11_c28 bl_28 br_28 wl_11 vdd gnd cell_6t
Xbit_r12_c28 bl_28 br_28 wl_12 vdd gnd cell_6t
Xbit_r13_c28 bl_28 br_28 wl_13 vdd gnd cell_6t
Xbit_r14_c28 bl_28 br_28 wl_14 vdd gnd cell_6t
Xbit_r15_c28 bl_28 br_28 wl_15 vdd gnd cell_6t
Xbit_r16_c28 bl_28 br_28 wl_16 vdd gnd cell_6t
Xbit_r17_c28 bl_28 br_28 wl_17 vdd gnd cell_6t
Xbit_r18_c28 bl_28 br_28 wl_18 vdd gnd cell_6t
Xbit_r19_c28 bl_28 br_28 wl_19 vdd gnd cell_6t
Xbit_r20_c28 bl_28 br_28 wl_20 vdd gnd cell_6t
Xbit_r21_c28 bl_28 br_28 wl_21 vdd gnd cell_6t
Xbit_r22_c28 bl_28 br_28 wl_22 vdd gnd cell_6t
Xbit_r23_c28 bl_28 br_28 wl_23 vdd gnd cell_6t
Xbit_r24_c28 bl_28 br_28 wl_24 vdd gnd cell_6t
Xbit_r25_c28 bl_28 br_28 wl_25 vdd gnd cell_6t
Xbit_r26_c28 bl_28 br_28 wl_26 vdd gnd cell_6t
Xbit_r27_c28 bl_28 br_28 wl_27 vdd gnd cell_6t
Xbit_r28_c28 bl_28 br_28 wl_28 vdd gnd cell_6t
Xbit_r29_c28 bl_28 br_28 wl_29 vdd gnd cell_6t
Xbit_r30_c28 bl_28 br_28 wl_30 vdd gnd cell_6t
Xbit_r31_c28 bl_28 br_28 wl_31 vdd gnd cell_6t
Xbit_r32_c28 bl_28 br_28 wl_32 vdd gnd cell_6t
Xbit_r33_c28 bl_28 br_28 wl_33 vdd gnd cell_6t
Xbit_r34_c28 bl_28 br_28 wl_34 vdd gnd cell_6t
Xbit_r35_c28 bl_28 br_28 wl_35 vdd gnd cell_6t
Xbit_r36_c28 bl_28 br_28 wl_36 vdd gnd cell_6t
Xbit_r37_c28 bl_28 br_28 wl_37 vdd gnd cell_6t
Xbit_r38_c28 bl_28 br_28 wl_38 vdd gnd cell_6t
Xbit_r39_c28 bl_28 br_28 wl_39 vdd gnd cell_6t
Xbit_r40_c28 bl_28 br_28 wl_40 vdd gnd cell_6t
Xbit_r41_c28 bl_28 br_28 wl_41 vdd gnd cell_6t
Xbit_r42_c28 bl_28 br_28 wl_42 vdd gnd cell_6t
Xbit_r43_c28 bl_28 br_28 wl_43 vdd gnd cell_6t
Xbit_r44_c28 bl_28 br_28 wl_44 vdd gnd cell_6t
Xbit_r45_c28 bl_28 br_28 wl_45 vdd gnd cell_6t
Xbit_r46_c28 bl_28 br_28 wl_46 vdd gnd cell_6t
Xbit_r47_c28 bl_28 br_28 wl_47 vdd gnd cell_6t
Xbit_r48_c28 bl_28 br_28 wl_48 vdd gnd cell_6t
Xbit_r49_c28 bl_28 br_28 wl_49 vdd gnd cell_6t
Xbit_r50_c28 bl_28 br_28 wl_50 vdd gnd cell_6t
Xbit_r51_c28 bl_28 br_28 wl_51 vdd gnd cell_6t
Xbit_r52_c28 bl_28 br_28 wl_52 vdd gnd cell_6t
Xbit_r53_c28 bl_28 br_28 wl_53 vdd gnd cell_6t
Xbit_r54_c28 bl_28 br_28 wl_54 vdd gnd cell_6t
Xbit_r55_c28 bl_28 br_28 wl_55 vdd gnd cell_6t
Xbit_r56_c28 bl_28 br_28 wl_56 vdd gnd cell_6t
Xbit_r57_c28 bl_28 br_28 wl_57 vdd gnd cell_6t
Xbit_r58_c28 bl_28 br_28 wl_58 vdd gnd cell_6t
Xbit_r59_c28 bl_28 br_28 wl_59 vdd gnd cell_6t
Xbit_r60_c28 bl_28 br_28 wl_60 vdd gnd cell_6t
Xbit_r61_c28 bl_28 br_28 wl_61 vdd gnd cell_6t
Xbit_r62_c28 bl_28 br_28 wl_62 vdd gnd cell_6t
Xbit_r63_c28 bl_28 br_28 wl_63 vdd gnd cell_6t
Xbit_r64_c28 bl_28 br_28 wl_64 vdd gnd cell_6t
Xbit_r65_c28 bl_28 br_28 wl_65 vdd gnd cell_6t
Xbit_r66_c28 bl_28 br_28 wl_66 vdd gnd cell_6t
Xbit_r67_c28 bl_28 br_28 wl_67 vdd gnd cell_6t
Xbit_r68_c28 bl_28 br_28 wl_68 vdd gnd cell_6t
Xbit_r69_c28 bl_28 br_28 wl_69 vdd gnd cell_6t
Xbit_r70_c28 bl_28 br_28 wl_70 vdd gnd cell_6t
Xbit_r71_c28 bl_28 br_28 wl_71 vdd gnd cell_6t
Xbit_r72_c28 bl_28 br_28 wl_72 vdd gnd cell_6t
Xbit_r73_c28 bl_28 br_28 wl_73 vdd gnd cell_6t
Xbit_r74_c28 bl_28 br_28 wl_74 vdd gnd cell_6t
Xbit_r75_c28 bl_28 br_28 wl_75 vdd gnd cell_6t
Xbit_r76_c28 bl_28 br_28 wl_76 vdd gnd cell_6t
Xbit_r77_c28 bl_28 br_28 wl_77 vdd gnd cell_6t
Xbit_r78_c28 bl_28 br_28 wl_78 vdd gnd cell_6t
Xbit_r79_c28 bl_28 br_28 wl_79 vdd gnd cell_6t
Xbit_r80_c28 bl_28 br_28 wl_80 vdd gnd cell_6t
Xbit_r81_c28 bl_28 br_28 wl_81 vdd gnd cell_6t
Xbit_r82_c28 bl_28 br_28 wl_82 vdd gnd cell_6t
Xbit_r83_c28 bl_28 br_28 wl_83 vdd gnd cell_6t
Xbit_r84_c28 bl_28 br_28 wl_84 vdd gnd cell_6t
Xbit_r85_c28 bl_28 br_28 wl_85 vdd gnd cell_6t
Xbit_r86_c28 bl_28 br_28 wl_86 vdd gnd cell_6t
Xbit_r87_c28 bl_28 br_28 wl_87 vdd gnd cell_6t
Xbit_r88_c28 bl_28 br_28 wl_88 vdd gnd cell_6t
Xbit_r89_c28 bl_28 br_28 wl_89 vdd gnd cell_6t
Xbit_r90_c28 bl_28 br_28 wl_90 vdd gnd cell_6t
Xbit_r91_c28 bl_28 br_28 wl_91 vdd gnd cell_6t
Xbit_r92_c28 bl_28 br_28 wl_92 vdd gnd cell_6t
Xbit_r93_c28 bl_28 br_28 wl_93 vdd gnd cell_6t
Xbit_r94_c28 bl_28 br_28 wl_94 vdd gnd cell_6t
Xbit_r95_c28 bl_28 br_28 wl_95 vdd gnd cell_6t
Xbit_r96_c28 bl_28 br_28 wl_96 vdd gnd cell_6t
Xbit_r97_c28 bl_28 br_28 wl_97 vdd gnd cell_6t
Xbit_r98_c28 bl_28 br_28 wl_98 vdd gnd cell_6t
Xbit_r99_c28 bl_28 br_28 wl_99 vdd gnd cell_6t
Xbit_r100_c28 bl_28 br_28 wl_100 vdd gnd cell_6t
Xbit_r101_c28 bl_28 br_28 wl_101 vdd gnd cell_6t
Xbit_r102_c28 bl_28 br_28 wl_102 vdd gnd cell_6t
Xbit_r103_c28 bl_28 br_28 wl_103 vdd gnd cell_6t
Xbit_r104_c28 bl_28 br_28 wl_104 vdd gnd cell_6t
Xbit_r105_c28 bl_28 br_28 wl_105 vdd gnd cell_6t
Xbit_r106_c28 bl_28 br_28 wl_106 vdd gnd cell_6t
Xbit_r107_c28 bl_28 br_28 wl_107 vdd gnd cell_6t
Xbit_r108_c28 bl_28 br_28 wl_108 vdd gnd cell_6t
Xbit_r109_c28 bl_28 br_28 wl_109 vdd gnd cell_6t
Xbit_r110_c28 bl_28 br_28 wl_110 vdd gnd cell_6t
Xbit_r111_c28 bl_28 br_28 wl_111 vdd gnd cell_6t
Xbit_r112_c28 bl_28 br_28 wl_112 vdd gnd cell_6t
Xbit_r113_c28 bl_28 br_28 wl_113 vdd gnd cell_6t
Xbit_r114_c28 bl_28 br_28 wl_114 vdd gnd cell_6t
Xbit_r115_c28 bl_28 br_28 wl_115 vdd gnd cell_6t
Xbit_r116_c28 bl_28 br_28 wl_116 vdd gnd cell_6t
Xbit_r117_c28 bl_28 br_28 wl_117 vdd gnd cell_6t
Xbit_r118_c28 bl_28 br_28 wl_118 vdd gnd cell_6t
Xbit_r119_c28 bl_28 br_28 wl_119 vdd gnd cell_6t
Xbit_r120_c28 bl_28 br_28 wl_120 vdd gnd cell_6t
Xbit_r121_c28 bl_28 br_28 wl_121 vdd gnd cell_6t
Xbit_r122_c28 bl_28 br_28 wl_122 vdd gnd cell_6t
Xbit_r123_c28 bl_28 br_28 wl_123 vdd gnd cell_6t
Xbit_r124_c28 bl_28 br_28 wl_124 vdd gnd cell_6t
Xbit_r125_c28 bl_28 br_28 wl_125 vdd gnd cell_6t
Xbit_r126_c28 bl_28 br_28 wl_126 vdd gnd cell_6t
Xbit_r127_c28 bl_28 br_28 wl_127 vdd gnd cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd cell_6t
Xbit_r1_c29 bl_29 br_29 wl_1 vdd gnd cell_6t
Xbit_r2_c29 bl_29 br_29 wl_2 vdd gnd cell_6t
Xbit_r3_c29 bl_29 br_29 wl_3 vdd gnd cell_6t
Xbit_r4_c29 bl_29 br_29 wl_4 vdd gnd cell_6t
Xbit_r5_c29 bl_29 br_29 wl_5 vdd gnd cell_6t
Xbit_r6_c29 bl_29 br_29 wl_6 vdd gnd cell_6t
Xbit_r7_c29 bl_29 br_29 wl_7 vdd gnd cell_6t
Xbit_r8_c29 bl_29 br_29 wl_8 vdd gnd cell_6t
Xbit_r9_c29 bl_29 br_29 wl_9 vdd gnd cell_6t
Xbit_r10_c29 bl_29 br_29 wl_10 vdd gnd cell_6t
Xbit_r11_c29 bl_29 br_29 wl_11 vdd gnd cell_6t
Xbit_r12_c29 bl_29 br_29 wl_12 vdd gnd cell_6t
Xbit_r13_c29 bl_29 br_29 wl_13 vdd gnd cell_6t
Xbit_r14_c29 bl_29 br_29 wl_14 vdd gnd cell_6t
Xbit_r15_c29 bl_29 br_29 wl_15 vdd gnd cell_6t
Xbit_r16_c29 bl_29 br_29 wl_16 vdd gnd cell_6t
Xbit_r17_c29 bl_29 br_29 wl_17 vdd gnd cell_6t
Xbit_r18_c29 bl_29 br_29 wl_18 vdd gnd cell_6t
Xbit_r19_c29 bl_29 br_29 wl_19 vdd gnd cell_6t
Xbit_r20_c29 bl_29 br_29 wl_20 vdd gnd cell_6t
Xbit_r21_c29 bl_29 br_29 wl_21 vdd gnd cell_6t
Xbit_r22_c29 bl_29 br_29 wl_22 vdd gnd cell_6t
Xbit_r23_c29 bl_29 br_29 wl_23 vdd gnd cell_6t
Xbit_r24_c29 bl_29 br_29 wl_24 vdd gnd cell_6t
Xbit_r25_c29 bl_29 br_29 wl_25 vdd gnd cell_6t
Xbit_r26_c29 bl_29 br_29 wl_26 vdd gnd cell_6t
Xbit_r27_c29 bl_29 br_29 wl_27 vdd gnd cell_6t
Xbit_r28_c29 bl_29 br_29 wl_28 vdd gnd cell_6t
Xbit_r29_c29 bl_29 br_29 wl_29 vdd gnd cell_6t
Xbit_r30_c29 bl_29 br_29 wl_30 vdd gnd cell_6t
Xbit_r31_c29 bl_29 br_29 wl_31 vdd gnd cell_6t
Xbit_r32_c29 bl_29 br_29 wl_32 vdd gnd cell_6t
Xbit_r33_c29 bl_29 br_29 wl_33 vdd gnd cell_6t
Xbit_r34_c29 bl_29 br_29 wl_34 vdd gnd cell_6t
Xbit_r35_c29 bl_29 br_29 wl_35 vdd gnd cell_6t
Xbit_r36_c29 bl_29 br_29 wl_36 vdd gnd cell_6t
Xbit_r37_c29 bl_29 br_29 wl_37 vdd gnd cell_6t
Xbit_r38_c29 bl_29 br_29 wl_38 vdd gnd cell_6t
Xbit_r39_c29 bl_29 br_29 wl_39 vdd gnd cell_6t
Xbit_r40_c29 bl_29 br_29 wl_40 vdd gnd cell_6t
Xbit_r41_c29 bl_29 br_29 wl_41 vdd gnd cell_6t
Xbit_r42_c29 bl_29 br_29 wl_42 vdd gnd cell_6t
Xbit_r43_c29 bl_29 br_29 wl_43 vdd gnd cell_6t
Xbit_r44_c29 bl_29 br_29 wl_44 vdd gnd cell_6t
Xbit_r45_c29 bl_29 br_29 wl_45 vdd gnd cell_6t
Xbit_r46_c29 bl_29 br_29 wl_46 vdd gnd cell_6t
Xbit_r47_c29 bl_29 br_29 wl_47 vdd gnd cell_6t
Xbit_r48_c29 bl_29 br_29 wl_48 vdd gnd cell_6t
Xbit_r49_c29 bl_29 br_29 wl_49 vdd gnd cell_6t
Xbit_r50_c29 bl_29 br_29 wl_50 vdd gnd cell_6t
Xbit_r51_c29 bl_29 br_29 wl_51 vdd gnd cell_6t
Xbit_r52_c29 bl_29 br_29 wl_52 vdd gnd cell_6t
Xbit_r53_c29 bl_29 br_29 wl_53 vdd gnd cell_6t
Xbit_r54_c29 bl_29 br_29 wl_54 vdd gnd cell_6t
Xbit_r55_c29 bl_29 br_29 wl_55 vdd gnd cell_6t
Xbit_r56_c29 bl_29 br_29 wl_56 vdd gnd cell_6t
Xbit_r57_c29 bl_29 br_29 wl_57 vdd gnd cell_6t
Xbit_r58_c29 bl_29 br_29 wl_58 vdd gnd cell_6t
Xbit_r59_c29 bl_29 br_29 wl_59 vdd gnd cell_6t
Xbit_r60_c29 bl_29 br_29 wl_60 vdd gnd cell_6t
Xbit_r61_c29 bl_29 br_29 wl_61 vdd gnd cell_6t
Xbit_r62_c29 bl_29 br_29 wl_62 vdd gnd cell_6t
Xbit_r63_c29 bl_29 br_29 wl_63 vdd gnd cell_6t
Xbit_r64_c29 bl_29 br_29 wl_64 vdd gnd cell_6t
Xbit_r65_c29 bl_29 br_29 wl_65 vdd gnd cell_6t
Xbit_r66_c29 bl_29 br_29 wl_66 vdd gnd cell_6t
Xbit_r67_c29 bl_29 br_29 wl_67 vdd gnd cell_6t
Xbit_r68_c29 bl_29 br_29 wl_68 vdd gnd cell_6t
Xbit_r69_c29 bl_29 br_29 wl_69 vdd gnd cell_6t
Xbit_r70_c29 bl_29 br_29 wl_70 vdd gnd cell_6t
Xbit_r71_c29 bl_29 br_29 wl_71 vdd gnd cell_6t
Xbit_r72_c29 bl_29 br_29 wl_72 vdd gnd cell_6t
Xbit_r73_c29 bl_29 br_29 wl_73 vdd gnd cell_6t
Xbit_r74_c29 bl_29 br_29 wl_74 vdd gnd cell_6t
Xbit_r75_c29 bl_29 br_29 wl_75 vdd gnd cell_6t
Xbit_r76_c29 bl_29 br_29 wl_76 vdd gnd cell_6t
Xbit_r77_c29 bl_29 br_29 wl_77 vdd gnd cell_6t
Xbit_r78_c29 bl_29 br_29 wl_78 vdd gnd cell_6t
Xbit_r79_c29 bl_29 br_29 wl_79 vdd gnd cell_6t
Xbit_r80_c29 bl_29 br_29 wl_80 vdd gnd cell_6t
Xbit_r81_c29 bl_29 br_29 wl_81 vdd gnd cell_6t
Xbit_r82_c29 bl_29 br_29 wl_82 vdd gnd cell_6t
Xbit_r83_c29 bl_29 br_29 wl_83 vdd gnd cell_6t
Xbit_r84_c29 bl_29 br_29 wl_84 vdd gnd cell_6t
Xbit_r85_c29 bl_29 br_29 wl_85 vdd gnd cell_6t
Xbit_r86_c29 bl_29 br_29 wl_86 vdd gnd cell_6t
Xbit_r87_c29 bl_29 br_29 wl_87 vdd gnd cell_6t
Xbit_r88_c29 bl_29 br_29 wl_88 vdd gnd cell_6t
Xbit_r89_c29 bl_29 br_29 wl_89 vdd gnd cell_6t
Xbit_r90_c29 bl_29 br_29 wl_90 vdd gnd cell_6t
Xbit_r91_c29 bl_29 br_29 wl_91 vdd gnd cell_6t
Xbit_r92_c29 bl_29 br_29 wl_92 vdd gnd cell_6t
Xbit_r93_c29 bl_29 br_29 wl_93 vdd gnd cell_6t
Xbit_r94_c29 bl_29 br_29 wl_94 vdd gnd cell_6t
Xbit_r95_c29 bl_29 br_29 wl_95 vdd gnd cell_6t
Xbit_r96_c29 bl_29 br_29 wl_96 vdd gnd cell_6t
Xbit_r97_c29 bl_29 br_29 wl_97 vdd gnd cell_6t
Xbit_r98_c29 bl_29 br_29 wl_98 vdd gnd cell_6t
Xbit_r99_c29 bl_29 br_29 wl_99 vdd gnd cell_6t
Xbit_r100_c29 bl_29 br_29 wl_100 vdd gnd cell_6t
Xbit_r101_c29 bl_29 br_29 wl_101 vdd gnd cell_6t
Xbit_r102_c29 bl_29 br_29 wl_102 vdd gnd cell_6t
Xbit_r103_c29 bl_29 br_29 wl_103 vdd gnd cell_6t
Xbit_r104_c29 bl_29 br_29 wl_104 vdd gnd cell_6t
Xbit_r105_c29 bl_29 br_29 wl_105 vdd gnd cell_6t
Xbit_r106_c29 bl_29 br_29 wl_106 vdd gnd cell_6t
Xbit_r107_c29 bl_29 br_29 wl_107 vdd gnd cell_6t
Xbit_r108_c29 bl_29 br_29 wl_108 vdd gnd cell_6t
Xbit_r109_c29 bl_29 br_29 wl_109 vdd gnd cell_6t
Xbit_r110_c29 bl_29 br_29 wl_110 vdd gnd cell_6t
Xbit_r111_c29 bl_29 br_29 wl_111 vdd gnd cell_6t
Xbit_r112_c29 bl_29 br_29 wl_112 vdd gnd cell_6t
Xbit_r113_c29 bl_29 br_29 wl_113 vdd gnd cell_6t
Xbit_r114_c29 bl_29 br_29 wl_114 vdd gnd cell_6t
Xbit_r115_c29 bl_29 br_29 wl_115 vdd gnd cell_6t
Xbit_r116_c29 bl_29 br_29 wl_116 vdd gnd cell_6t
Xbit_r117_c29 bl_29 br_29 wl_117 vdd gnd cell_6t
Xbit_r118_c29 bl_29 br_29 wl_118 vdd gnd cell_6t
Xbit_r119_c29 bl_29 br_29 wl_119 vdd gnd cell_6t
Xbit_r120_c29 bl_29 br_29 wl_120 vdd gnd cell_6t
Xbit_r121_c29 bl_29 br_29 wl_121 vdd gnd cell_6t
Xbit_r122_c29 bl_29 br_29 wl_122 vdd gnd cell_6t
Xbit_r123_c29 bl_29 br_29 wl_123 vdd gnd cell_6t
Xbit_r124_c29 bl_29 br_29 wl_124 vdd gnd cell_6t
Xbit_r125_c29 bl_29 br_29 wl_125 vdd gnd cell_6t
Xbit_r126_c29 bl_29 br_29 wl_126 vdd gnd cell_6t
Xbit_r127_c29 bl_29 br_29 wl_127 vdd gnd cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd cell_6t
Xbit_r1_c30 bl_30 br_30 wl_1 vdd gnd cell_6t
Xbit_r2_c30 bl_30 br_30 wl_2 vdd gnd cell_6t
Xbit_r3_c30 bl_30 br_30 wl_3 vdd gnd cell_6t
Xbit_r4_c30 bl_30 br_30 wl_4 vdd gnd cell_6t
Xbit_r5_c30 bl_30 br_30 wl_5 vdd gnd cell_6t
Xbit_r6_c30 bl_30 br_30 wl_6 vdd gnd cell_6t
Xbit_r7_c30 bl_30 br_30 wl_7 vdd gnd cell_6t
Xbit_r8_c30 bl_30 br_30 wl_8 vdd gnd cell_6t
Xbit_r9_c30 bl_30 br_30 wl_9 vdd gnd cell_6t
Xbit_r10_c30 bl_30 br_30 wl_10 vdd gnd cell_6t
Xbit_r11_c30 bl_30 br_30 wl_11 vdd gnd cell_6t
Xbit_r12_c30 bl_30 br_30 wl_12 vdd gnd cell_6t
Xbit_r13_c30 bl_30 br_30 wl_13 vdd gnd cell_6t
Xbit_r14_c30 bl_30 br_30 wl_14 vdd gnd cell_6t
Xbit_r15_c30 bl_30 br_30 wl_15 vdd gnd cell_6t
Xbit_r16_c30 bl_30 br_30 wl_16 vdd gnd cell_6t
Xbit_r17_c30 bl_30 br_30 wl_17 vdd gnd cell_6t
Xbit_r18_c30 bl_30 br_30 wl_18 vdd gnd cell_6t
Xbit_r19_c30 bl_30 br_30 wl_19 vdd gnd cell_6t
Xbit_r20_c30 bl_30 br_30 wl_20 vdd gnd cell_6t
Xbit_r21_c30 bl_30 br_30 wl_21 vdd gnd cell_6t
Xbit_r22_c30 bl_30 br_30 wl_22 vdd gnd cell_6t
Xbit_r23_c30 bl_30 br_30 wl_23 vdd gnd cell_6t
Xbit_r24_c30 bl_30 br_30 wl_24 vdd gnd cell_6t
Xbit_r25_c30 bl_30 br_30 wl_25 vdd gnd cell_6t
Xbit_r26_c30 bl_30 br_30 wl_26 vdd gnd cell_6t
Xbit_r27_c30 bl_30 br_30 wl_27 vdd gnd cell_6t
Xbit_r28_c30 bl_30 br_30 wl_28 vdd gnd cell_6t
Xbit_r29_c30 bl_30 br_30 wl_29 vdd gnd cell_6t
Xbit_r30_c30 bl_30 br_30 wl_30 vdd gnd cell_6t
Xbit_r31_c30 bl_30 br_30 wl_31 vdd gnd cell_6t
Xbit_r32_c30 bl_30 br_30 wl_32 vdd gnd cell_6t
Xbit_r33_c30 bl_30 br_30 wl_33 vdd gnd cell_6t
Xbit_r34_c30 bl_30 br_30 wl_34 vdd gnd cell_6t
Xbit_r35_c30 bl_30 br_30 wl_35 vdd gnd cell_6t
Xbit_r36_c30 bl_30 br_30 wl_36 vdd gnd cell_6t
Xbit_r37_c30 bl_30 br_30 wl_37 vdd gnd cell_6t
Xbit_r38_c30 bl_30 br_30 wl_38 vdd gnd cell_6t
Xbit_r39_c30 bl_30 br_30 wl_39 vdd gnd cell_6t
Xbit_r40_c30 bl_30 br_30 wl_40 vdd gnd cell_6t
Xbit_r41_c30 bl_30 br_30 wl_41 vdd gnd cell_6t
Xbit_r42_c30 bl_30 br_30 wl_42 vdd gnd cell_6t
Xbit_r43_c30 bl_30 br_30 wl_43 vdd gnd cell_6t
Xbit_r44_c30 bl_30 br_30 wl_44 vdd gnd cell_6t
Xbit_r45_c30 bl_30 br_30 wl_45 vdd gnd cell_6t
Xbit_r46_c30 bl_30 br_30 wl_46 vdd gnd cell_6t
Xbit_r47_c30 bl_30 br_30 wl_47 vdd gnd cell_6t
Xbit_r48_c30 bl_30 br_30 wl_48 vdd gnd cell_6t
Xbit_r49_c30 bl_30 br_30 wl_49 vdd gnd cell_6t
Xbit_r50_c30 bl_30 br_30 wl_50 vdd gnd cell_6t
Xbit_r51_c30 bl_30 br_30 wl_51 vdd gnd cell_6t
Xbit_r52_c30 bl_30 br_30 wl_52 vdd gnd cell_6t
Xbit_r53_c30 bl_30 br_30 wl_53 vdd gnd cell_6t
Xbit_r54_c30 bl_30 br_30 wl_54 vdd gnd cell_6t
Xbit_r55_c30 bl_30 br_30 wl_55 vdd gnd cell_6t
Xbit_r56_c30 bl_30 br_30 wl_56 vdd gnd cell_6t
Xbit_r57_c30 bl_30 br_30 wl_57 vdd gnd cell_6t
Xbit_r58_c30 bl_30 br_30 wl_58 vdd gnd cell_6t
Xbit_r59_c30 bl_30 br_30 wl_59 vdd gnd cell_6t
Xbit_r60_c30 bl_30 br_30 wl_60 vdd gnd cell_6t
Xbit_r61_c30 bl_30 br_30 wl_61 vdd gnd cell_6t
Xbit_r62_c30 bl_30 br_30 wl_62 vdd gnd cell_6t
Xbit_r63_c30 bl_30 br_30 wl_63 vdd gnd cell_6t
Xbit_r64_c30 bl_30 br_30 wl_64 vdd gnd cell_6t
Xbit_r65_c30 bl_30 br_30 wl_65 vdd gnd cell_6t
Xbit_r66_c30 bl_30 br_30 wl_66 vdd gnd cell_6t
Xbit_r67_c30 bl_30 br_30 wl_67 vdd gnd cell_6t
Xbit_r68_c30 bl_30 br_30 wl_68 vdd gnd cell_6t
Xbit_r69_c30 bl_30 br_30 wl_69 vdd gnd cell_6t
Xbit_r70_c30 bl_30 br_30 wl_70 vdd gnd cell_6t
Xbit_r71_c30 bl_30 br_30 wl_71 vdd gnd cell_6t
Xbit_r72_c30 bl_30 br_30 wl_72 vdd gnd cell_6t
Xbit_r73_c30 bl_30 br_30 wl_73 vdd gnd cell_6t
Xbit_r74_c30 bl_30 br_30 wl_74 vdd gnd cell_6t
Xbit_r75_c30 bl_30 br_30 wl_75 vdd gnd cell_6t
Xbit_r76_c30 bl_30 br_30 wl_76 vdd gnd cell_6t
Xbit_r77_c30 bl_30 br_30 wl_77 vdd gnd cell_6t
Xbit_r78_c30 bl_30 br_30 wl_78 vdd gnd cell_6t
Xbit_r79_c30 bl_30 br_30 wl_79 vdd gnd cell_6t
Xbit_r80_c30 bl_30 br_30 wl_80 vdd gnd cell_6t
Xbit_r81_c30 bl_30 br_30 wl_81 vdd gnd cell_6t
Xbit_r82_c30 bl_30 br_30 wl_82 vdd gnd cell_6t
Xbit_r83_c30 bl_30 br_30 wl_83 vdd gnd cell_6t
Xbit_r84_c30 bl_30 br_30 wl_84 vdd gnd cell_6t
Xbit_r85_c30 bl_30 br_30 wl_85 vdd gnd cell_6t
Xbit_r86_c30 bl_30 br_30 wl_86 vdd gnd cell_6t
Xbit_r87_c30 bl_30 br_30 wl_87 vdd gnd cell_6t
Xbit_r88_c30 bl_30 br_30 wl_88 vdd gnd cell_6t
Xbit_r89_c30 bl_30 br_30 wl_89 vdd gnd cell_6t
Xbit_r90_c30 bl_30 br_30 wl_90 vdd gnd cell_6t
Xbit_r91_c30 bl_30 br_30 wl_91 vdd gnd cell_6t
Xbit_r92_c30 bl_30 br_30 wl_92 vdd gnd cell_6t
Xbit_r93_c30 bl_30 br_30 wl_93 vdd gnd cell_6t
Xbit_r94_c30 bl_30 br_30 wl_94 vdd gnd cell_6t
Xbit_r95_c30 bl_30 br_30 wl_95 vdd gnd cell_6t
Xbit_r96_c30 bl_30 br_30 wl_96 vdd gnd cell_6t
Xbit_r97_c30 bl_30 br_30 wl_97 vdd gnd cell_6t
Xbit_r98_c30 bl_30 br_30 wl_98 vdd gnd cell_6t
Xbit_r99_c30 bl_30 br_30 wl_99 vdd gnd cell_6t
Xbit_r100_c30 bl_30 br_30 wl_100 vdd gnd cell_6t
Xbit_r101_c30 bl_30 br_30 wl_101 vdd gnd cell_6t
Xbit_r102_c30 bl_30 br_30 wl_102 vdd gnd cell_6t
Xbit_r103_c30 bl_30 br_30 wl_103 vdd gnd cell_6t
Xbit_r104_c30 bl_30 br_30 wl_104 vdd gnd cell_6t
Xbit_r105_c30 bl_30 br_30 wl_105 vdd gnd cell_6t
Xbit_r106_c30 bl_30 br_30 wl_106 vdd gnd cell_6t
Xbit_r107_c30 bl_30 br_30 wl_107 vdd gnd cell_6t
Xbit_r108_c30 bl_30 br_30 wl_108 vdd gnd cell_6t
Xbit_r109_c30 bl_30 br_30 wl_109 vdd gnd cell_6t
Xbit_r110_c30 bl_30 br_30 wl_110 vdd gnd cell_6t
Xbit_r111_c30 bl_30 br_30 wl_111 vdd gnd cell_6t
Xbit_r112_c30 bl_30 br_30 wl_112 vdd gnd cell_6t
Xbit_r113_c30 bl_30 br_30 wl_113 vdd gnd cell_6t
Xbit_r114_c30 bl_30 br_30 wl_114 vdd gnd cell_6t
Xbit_r115_c30 bl_30 br_30 wl_115 vdd gnd cell_6t
Xbit_r116_c30 bl_30 br_30 wl_116 vdd gnd cell_6t
Xbit_r117_c30 bl_30 br_30 wl_117 vdd gnd cell_6t
Xbit_r118_c30 bl_30 br_30 wl_118 vdd gnd cell_6t
Xbit_r119_c30 bl_30 br_30 wl_119 vdd gnd cell_6t
Xbit_r120_c30 bl_30 br_30 wl_120 vdd gnd cell_6t
Xbit_r121_c30 bl_30 br_30 wl_121 vdd gnd cell_6t
Xbit_r122_c30 bl_30 br_30 wl_122 vdd gnd cell_6t
Xbit_r123_c30 bl_30 br_30 wl_123 vdd gnd cell_6t
Xbit_r124_c30 bl_30 br_30 wl_124 vdd gnd cell_6t
Xbit_r125_c30 bl_30 br_30 wl_125 vdd gnd cell_6t
Xbit_r126_c30 bl_30 br_30 wl_126 vdd gnd cell_6t
Xbit_r127_c30 bl_30 br_30 wl_127 vdd gnd cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd cell_6t
Xbit_r1_c31 bl_31 br_31 wl_1 vdd gnd cell_6t
Xbit_r2_c31 bl_31 br_31 wl_2 vdd gnd cell_6t
Xbit_r3_c31 bl_31 br_31 wl_3 vdd gnd cell_6t
Xbit_r4_c31 bl_31 br_31 wl_4 vdd gnd cell_6t
Xbit_r5_c31 bl_31 br_31 wl_5 vdd gnd cell_6t
Xbit_r6_c31 bl_31 br_31 wl_6 vdd gnd cell_6t
Xbit_r7_c31 bl_31 br_31 wl_7 vdd gnd cell_6t
Xbit_r8_c31 bl_31 br_31 wl_8 vdd gnd cell_6t
Xbit_r9_c31 bl_31 br_31 wl_9 vdd gnd cell_6t
Xbit_r10_c31 bl_31 br_31 wl_10 vdd gnd cell_6t
Xbit_r11_c31 bl_31 br_31 wl_11 vdd gnd cell_6t
Xbit_r12_c31 bl_31 br_31 wl_12 vdd gnd cell_6t
Xbit_r13_c31 bl_31 br_31 wl_13 vdd gnd cell_6t
Xbit_r14_c31 bl_31 br_31 wl_14 vdd gnd cell_6t
Xbit_r15_c31 bl_31 br_31 wl_15 vdd gnd cell_6t
Xbit_r16_c31 bl_31 br_31 wl_16 vdd gnd cell_6t
Xbit_r17_c31 bl_31 br_31 wl_17 vdd gnd cell_6t
Xbit_r18_c31 bl_31 br_31 wl_18 vdd gnd cell_6t
Xbit_r19_c31 bl_31 br_31 wl_19 vdd gnd cell_6t
Xbit_r20_c31 bl_31 br_31 wl_20 vdd gnd cell_6t
Xbit_r21_c31 bl_31 br_31 wl_21 vdd gnd cell_6t
Xbit_r22_c31 bl_31 br_31 wl_22 vdd gnd cell_6t
Xbit_r23_c31 bl_31 br_31 wl_23 vdd gnd cell_6t
Xbit_r24_c31 bl_31 br_31 wl_24 vdd gnd cell_6t
Xbit_r25_c31 bl_31 br_31 wl_25 vdd gnd cell_6t
Xbit_r26_c31 bl_31 br_31 wl_26 vdd gnd cell_6t
Xbit_r27_c31 bl_31 br_31 wl_27 vdd gnd cell_6t
Xbit_r28_c31 bl_31 br_31 wl_28 vdd gnd cell_6t
Xbit_r29_c31 bl_31 br_31 wl_29 vdd gnd cell_6t
Xbit_r30_c31 bl_31 br_31 wl_30 vdd gnd cell_6t
Xbit_r31_c31 bl_31 br_31 wl_31 vdd gnd cell_6t
Xbit_r32_c31 bl_31 br_31 wl_32 vdd gnd cell_6t
Xbit_r33_c31 bl_31 br_31 wl_33 vdd gnd cell_6t
Xbit_r34_c31 bl_31 br_31 wl_34 vdd gnd cell_6t
Xbit_r35_c31 bl_31 br_31 wl_35 vdd gnd cell_6t
Xbit_r36_c31 bl_31 br_31 wl_36 vdd gnd cell_6t
Xbit_r37_c31 bl_31 br_31 wl_37 vdd gnd cell_6t
Xbit_r38_c31 bl_31 br_31 wl_38 vdd gnd cell_6t
Xbit_r39_c31 bl_31 br_31 wl_39 vdd gnd cell_6t
Xbit_r40_c31 bl_31 br_31 wl_40 vdd gnd cell_6t
Xbit_r41_c31 bl_31 br_31 wl_41 vdd gnd cell_6t
Xbit_r42_c31 bl_31 br_31 wl_42 vdd gnd cell_6t
Xbit_r43_c31 bl_31 br_31 wl_43 vdd gnd cell_6t
Xbit_r44_c31 bl_31 br_31 wl_44 vdd gnd cell_6t
Xbit_r45_c31 bl_31 br_31 wl_45 vdd gnd cell_6t
Xbit_r46_c31 bl_31 br_31 wl_46 vdd gnd cell_6t
Xbit_r47_c31 bl_31 br_31 wl_47 vdd gnd cell_6t
Xbit_r48_c31 bl_31 br_31 wl_48 vdd gnd cell_6t
Xbit_r49_c31 bl_31 br_31 wl_49 vdd gnd cell_6t
Xbit_r50_c31 bl_31 br_31 wl_50 vdd gnd cell_6t
Xbit_r51_c31 bl_31 br_31 wl_51 vdd gnd cell_6t
Xbit_r52_c31 bl_31 br_31 wl_52 vdd gnd cell_6t
Xbit_r53_c31 bl_31 br_31 wl_53 vdd gnd cell_6t
Xbit_r54_c31 bl_31 br_31 wl_54 vdd gnd cell_6t
Xbit_r55_c31 bl_31 br_31 wl_55 vdd gnd cell_6t
Xbit_r56_c31 bl_31 br_31 wl_56 vdd gnd cell_6t
Xbit_r57_c31 bl_31 br_31 wl_57 vdd gnd cell_6t
Xbit_r58_c31 bl_31 br_31 wl_58 vdd gnd cell_6t
Xbit_r59_c31 bl_31 br_31 wl_59 vdd gnd cell_6t
Xbit_r60_c31 bl_31 br_31 wl_60 vdd gnd cell_6t
Xbit_r61_c31 bl_31 br_31 wl_61 vdd gnd cell_6t
Xbit_r62_c31 bl_31 br_31 wl_62 vdd gnd cell_6t
Xbit_r63_c31 bl_31 br_31 wl_63 vdd gnd cell_6t
Xbit_r64_c31 bl_31 br_31 wl_64 vdd gnd cell_6t
Xbit_r65_c31 bl_31 br_31 wl_65 vdd gnd cell_6t
Xbit_r66_c31 bl_31 br_31 wl_66 vdd gnd cell_6t
Xbit_r67_c31 bl_31 br_31 wl_67 vdd gnd cell_6t
Xbit_r68_c31 bl_31 br_31 wl_68 vdd gnd cell_6t
Xbit_r69_c31 bl_31 br_31 wl_69 vdd gnd cell_6t
Xbit_r70_c31 bl_31 br_31 wl_70 vdd gnd cell_6t
Xbit_r71_c31 bl_31 br_31 wl_71 vdd gnd cell_6t
Xbit_r72_c31 bl_31 br_31 wl_72 vdd gnd cell_6t
Xbit_r73_c31 bl_31 br_31 wl_73 vdd gnd cell_6t
Xbit_r74_c31 bl_31 br_31 wl_74 vdd gnd cell_6t
Xbit_r75_c31 bl_31 br_31 wl_75 vdd gnd cell_6t
Xbit_r76_c31 bl_31 br_31 wl_76 vdd gnd cell_6t
Xbit_r77_c31 bl_31 br_31 wl_77 vdd gnd cell_6t
Xbit_r78_c31 bl_31 br_31 wl_78 vdd gnd cell_6t
Xbit_r79_c31 bl_31 br_31 wl_79 vdd gnd cell_6t
Xbit_r80_c31 bl_31 br_31 wl_80 vdd gnd cell_6t
Xbit_r81_c31 bl_31 br_31 wl_81 vdd gnd cell_6t
Xbit_r82_c31 bl_31 br_31 wl_82 vdd gnd cell_6t
Xbit_r83_c31 bl_31 br_31 wl_83 vdd gnd cell_6t
Xbit_r84_c31 bl_31 br_31 wl_84 vdd gnd cell_6t
Xbit_r85_c31 bl_31 br_31 wl_85 vdd gnd cell_6t
Xbit_r86_c31 bl_31 br_31 wl_86 vdd gnd cell_6t
Xbit_r87_c31 bl_31 br_31 wl_87 vdd gnd cell_6t
Xbit_r88_c31 bl_31 br_31 wl_88 vdd gnd cell_6t
Xbit_r89_c31 bl_31 br_31 wl_89 vdd gnd cell_6t
Xbit_r90_c31 bl_31 br_31 wl_90 vdd gnd cell_6t
Xbit_r91_c31 bl_31 br_31 wl_91 vdd gnd cell_6t
Xbit_r92_c31 bl_31 br_31 wl_92 vdd gnd cell_6t
Xbit_r93_c31 bl_31 br_31 wl_93 vdd gnd cell_6t
Xbit_r94_c31 bl_31 br_31 wl_94 vdd gnd cell_6t
Xbit_r95_c31 bl_31 br_31 wl_95 vdd gnd cell_6t
Xbit_r96_c31 bl_31 br_31 wl_96 vdd gnd cell_6t
Xbit_r97_c31 bl_31 br_31 wl_97 vdd gnd cell_6t
Xbit_r98_c31 bl_31 br_31 wl_98 vdd gnd cell_6t
Xbit_r99_c31 bl_31 br_31 wl_99 vdd gnd cell_6t
Xbit_r100_c31 bl_31 br_31 wl_100 vdd gnd cell_6t
Xbit_r101_c31 bl_31 br_31 wl_101 vdd gnd cell_6t
Xbit_r102_c31 bl_31 br_31 wl_102 vdd gnd cell_6t
Xbit_r103_c31 bl_31 br_31 wl_103 vdd gnd cell_6t
Xbit_r104_c31 bl_31 br_31 wl_104 vdd gnd cell_6t
Xbit_r105_c31 bl_31 br_31 wl_105 vdd gnd cell_6t
Xbit_r106_c31 bl_31 br_31 wl_106 vdd gnd cell_6t
Xbit_r107_c31 bl_31 br_31 wl_107 vdd gnd cell_6t
Xbit_r108_c31 bl_31 br_31 wl_108 vdd gnd cell_6t
Xbit_r109_c31 bl_31 br_31 wl_109 vdd gnd cell_6t
Xbit_r110_c31 bl_31 br_31 wl_110 vdd gnd cell_6t
Xbit_r111_c31 bl_31 br_31 wl_111 vdd gnd cell_6t
Xbit_r112_c31 bl_31 br_31 wl_112 vdd gnd cell_6t
Xbit_r113_c31 bl_31 br_31 wl_113 vdd gnd cell_6t
Xbit_r114_c31 bl_31 br_31 wl_114 vdd gnd cell_6t
Xbit_r115_c31 bl_31 br_31 wl_115 vdd gnd cell_6t
Xbit_r116_c31 bl_31 br_31 wl_116 vdd gnd cell_6t
Xbit_r117_c31 bl_31 br_31 wl_117 vdd gnd cell_6t
Xbit_r118_c31 bl_31 br_31 wl_118 vdd gnd cell_6t
Xbit_r119_c31 bl_31 br_31 wl_119 vdd gnd cell_6t
Xbit_r120_c31 bl_31 br_31 wl_120 vdd gnd cell_6t
Xbit_r121_c31 bl_31 br_31 wl_121 vdd gnd cell_6t
Xbit_r122_c31 bl_31 br_31 wl_122 vdd gnd cell_6t
Xbit_r123_c31 bl_31 br_31 wl_123 vdd gnd cell_6t
Xbit_r124_c31 bl_31 br_31 wl_124 vdd gnd cell_6t
Xbit_r125_c31 bl_31 br_31 wl_125 vdd gnd cell_6t
Xbit_r126_c31 bl_31 br_31 wl_126 vdd gnd cell_6t
Xbit_r127_c31 bl_31 br_31 wl_127 vdd gnd cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd cell_6t
Xbit_r1_c32 bl_32 br_32 wl_1 vdd gnd cell_6t
Xbit_r2_c32 bl_32 br_32 wl_2 vdd gnd cell_6t
Xbit_r3_c32 bl_32 br_32 wl_3 vdd gnd cell_6t
Xbit_r4_c32 bl_32 br_32 wl_4 vdd gnd cell_6t
Xbit_r5_c32 bl_32 br_32 wl_5 vdd gnd cell_6t
Xbit_r6_c32 bl_32 br_32 wl_6 vdd gnd cell_6t
Xbit_r7_c32 bl_32 br_32 wl_7 vdd gnd cell_6t
Xbit_r8_c32 bl_32 br_32 wl_8 vdd gnd cell_6t
Xbit_r9_c32 bl_32 br_32 wl_9 vdd gnd cell_6t
Xbit_r10_c32 bl_32 br_32 wl_10 vdd gnd cell_6t
Xbit_r11_c32 bl_32 br_32 wl_11 vdd gnd cell_6t
Xbit_r12_c32 bl_32 br_32 wl_12 vdd gnd cell_6t
Xbit_r13_c32 bl_32 br_32 wl_13 vdd gnd cell_6t
Xbit_r14_c32 bl_32 br_32 wl_14 vdd gnd cell_6t
Xbit_r15_c32 bl_32 br_32 wl_15 vdd gnd cell_6t
Xbit_r16_c32 bl_32 br_32 wl_16 vdd gnd cell_6t
Xbit_r17_c32 bl_32 br_32 wl_17 vdd gnd cell_6t
Xbit_r18_c32 bl_32 br_32 wl_18 vdd gnd cell_6t
Xbit_r19_c32 bl_32 br_32 wl_19 vdd gnd cell_6t
Xbit_r20_c32 bl_32 br_32 wl_20 vdd gnd cell_6t
Xbit_r21_c32 bl_32 br_32 wl_21 vdd gnd cell_6t
Xbit_r22_c32 bl_32 br_32 wl_22 vdd gnd cell_6t
Xbit_r23_c32 bl_32 br_32 wl_23 vdd gnd cell_6t
Xbit_r24_c32 bl_32 br_32 wl_24 vdd gnd cell_6t
Xbit_r25_c32 bl_32 br_32 wl_25 vdd gnd cell_6t
Xbit_r26_c32 bl_32 br_32 wl_26 vdd gnd cell_6t
Xbit_r27_c32 bl_32 br_32 wl_27 vdd gnd cell_6t
Xbit_r28_c32 bl_32 br_32 wl_28 vdd gnd cell_6t
Xbit_r29_c32 bl_32 br_32 wl_29 vdd gnd cell_6t
Xbit_r30_c32 bl_32 br_32 wl_30 vdd gnd cell_6t
Xbit_r31_c32 bl_32 br_32 wl_31 vdd gnd cell_6t
Xbit_r32_c32 bl_32 br_32 wl_32 vdd gnd cell_6t
Xbit_r33_c32 bl_32 br_32 wl_33 vdd gnd cell_6t
Xbit_r34_c32 bl_32 br_32 wl_34 vdd gnd cell_6t
Xbit_r35_c32 bl_32 br_32 wl_35 vdd gnd cell_6t
Xbit_r36_c32 bl_32 br_32 wl_36 vdd gnd cell_6t
Xbit_r37_c32 bl_32 br_32 wl_37 vdd gnd cell_6t
Xbit_r38_c32 bl_32 br_32 wl_38 vdd gnd cell_6t
Xbit_r39_c32 bl_32 br_32 wl_39 vdd gnd cell_6t
Xbit_r40_c32 bl_32 br_32 wl_40 vdd gnd cell_6t
Xbit_r41_c32 bl_32 br_32 wl_41 vdd gnd cell_6t
Xbit_r42_c32 bl_32 br_32 wl_42 vdd gnd cell_6t
Xbit_r43_c32 bl_32 br_32 wl_43 vdd gnd cell_6t
Xbit_r44_c32 bl_32 br_32 wl_44 vdd gnd cell_6t
Xbit_r45_c32 bl_32 br_32 wl_45 vdd gnd cell_6t
Xbit_r46_c32 bl_32 br_32 wl_46 vdd gnd cell_6t
Xbit_r47_c32 bl_32 br_32 wl_47 vdd gnd cell_6t
Xbit_r48_c32 bl_32 br_32 wl_48 vdd gnd cell_6t
Xbit_r49_c32 bl_32 br_32 wl_49 vdd gnd cell_6t
Xbit_r50_c32 bl_32 br_32 wl_50 vdd gnd cell_6t
Xbit_r51_c32 bl_32 br_32 wl_51 vdd gnd cell_6t
Xbit_r52_c32 bl_32 br_32 wl_52 vdd gnd cell_6t
Xbit_r53_c32 bl_32 br_32 wl_53 vdd gnd cell_6t
Xbit_r54_c32 bl_32 br_32 wl_54 vdd gnd cell_6t
Xbit_r55_c32 bl_32 br_32 wl_55 vdd gnd cell_6t
Xbit_r56_c32 bl_32 br_32 wl_56 vdd gnd cell_6t
Xbit_r57_c32 bl_32 br_32 wl_57 vdd gnd cell_6t
Xbit_r58_c32 bl_32 br_32 wl_58 vdd gnd cell_6t
Xbit_r59_c32 bl_32 br_32 wl_59 vdd gnd cell_6t
Xbit_r60_c32 bl_32 br_32 wl_60 vdd gnd cell_6t
Xbit_r61_c32 bl_32 br_32 wl_61 vdd gnd cell_6t
Xbit_r62_c32 bl_32 br_32 wl_62 vdd gnd cell_6t
Xbit_r63_c32 bl_32 br_32 wl_63 vdd gnd cell_6t
Xbit_r64_c32 bl_32 br_32 wl_64 vdd gnd cell_6t
Xbit_r65_c32 bl_32 br_32 wl_65 vdd gnd cell_6t
Xbit_r66_c32 bl_32 br_32 wl_66 vdd gnd cell_6t
Xbit_r67_c32 bl_32 br_32 wl_67 vdd gnd cell_6t
Xbit_r68_c32 bl_32 br_32 wl_68 vdd gnd cell_6t
Xbit_r69_c32 bl_32 br_32 wl_69 vdd gnd cell_6t
Xbit_r70_c32 bl_32 br_32 wl_70 vdd gnd cell_6t
Xbit_r71_c32 bl_32 br_32 wl_71 vdd gnd cell_6t
Xbit_r72_c32 bl_32 br_32 wl_72 vdd gnd cell_6t
Xbit_r73_c32 bl_32 br_32 wl_73 vdd gnd cell_6t
Xbit_r74_c32 bl_32 br_32 wl_74 vdd gnd cell_6t
Xbit_r75_c32 bl_32 br_32 wl_75 vdd gnd cell_6t
Xbit_r76_c32 bl_32 br_32 wl_76 vdd gnd cell_6t
Xbit_r77_c32 bl_32 br_32 wl_77 vdd gnd cell_6t
Xbit_r78_c32 bl_32 br_32 wl_78 vdd gnd cell_6t
Xbit_r79_c32 bl_32 br_32 wl_79 vdd gnd cell_6t
Xbit_r80_c32 bl_32 br_32 wl_80 vdd gnd cell_6t
Xbit_r81_c32 bl_32 br_32 wl_81 vdd gnd cell_6t
Xbit_r82_c32 bl_32 br_32 wl_82 vdd gnd cell_6t
Xbit_r83_c32 bl_32 br_32 wl_83 vdd gnd cell_6t
Xbit_r84_c32 bl_32 br_32 wl_84 vdd gnd cell_6t
Xbit_r85_c32 bl_32 br_32 wl_85 vdd gnd cell_6t
Xbit_r86_c32 bl_32 br_32 wl_86 vdd gnd cell_6t
Xbit_r87_c32 bl_32 br_32 wl_87 vdd gnd cell_6t
Xbit_r88_c32 bl_32 br_32 wl_88 vdd gnd cell_6t
Xbit_r89_c32 bl_32 br_32 wl_89 vdd gnd cell_6t
Xbit_r90_c32 bl_32 br_32 wl_90 vdd gnd cell_6t
Xbit_r91_c32 bl_32 br_32 wl_91 vdd gnd cell_6t
Xbit_r92_c32 bl_32 br_32 wl_92 vdd gnd cell_6t
Xbit_r93_c32 bl_32 br_32 wl_93 vdd gnd cell_6t
Xbit_r94_c32 bl_32 br_32 wl_94 vdd gnd cell_6t
Xbit_r95_c32 bl_32 br_32 wl_95 vdd gnd cell_6t
Xbit_r96_c32 bl_32 br_32 wl_96 vdd gnd cell_6t
Xbit_r97_c32 bl_32 br_32 wl_97 vdd gnd cell_6t
Xbit_r98_c32 bl_32 br_32 wl_98 vdd gnd cell_6t
Xbit_r99_c32 bl_32 br_32 wl_99 vdd gnd cell_6t
Xbit_r100_c32 bl_32 br_32 wl_100 vdd gnd cell_6t
Xbit_r101_c32 bl_32 br_32 wl_101 vdd gnd cell_6t
Xbit_r102_c32 bl_32 br_32 wl_102 vdd gnd cell_6t
Xbit_r103_c32 bl_32 br_32 wl_103 vdd gnd cell_6t
Xbit_r104_c32 bl_32 br_32 wl_104 vdd gnd cell_6t
Xbit_r105_c32 bl_32 br_32 wl_105 vdd gnd cell_6t
Xbit_r106_c32 bl_32 br_32 wl_106 vdd gnd cell_6t
Xbit_r107_c32 bl_32 br_32 wl_107 vdd gnd cell_6t
Xbit_r108_c32 bl_32 br_32 wl_108 vdd gnd cell_6t
Xbit_r109_c32 bl_32 br_32 wl_109 vdd gnd cell_6t
Xbit_r110_c32 bl_32 br_32 wl_110 vdd gnd cell_6t
Xbit_r111_c32 bl_32 br_32 wl_111 vdd gnd cell_6t
Xbit_r112_c32 bl_32 br_32 wl_112 vdd gnd cell_6t
Xbit_r113_c32 bl_32 br_32 wl_113 vdd gnd cell_6t
Xbit_r114_c32 bl_32 br_32 wl_114 vdd gnd cell_6t
Xbit_r115_c32 bl_32 br_32 wl_115 vdd gnd cell_6t
Xbit_r116_c32 bl_32 br_32 wl_116 vdd gnd cell_6t
Xbit_r117_c32 bl_32 br_32 wl_117 vdd gnd cell_6t
Xbit_r118_c32 bl_32 br_32 wl_118 vdd gnd cell_6t
Xbit_r119_c32 bl_32 br_32 wl_119 vdd gnd cell_6t
Xbit_r120_c32 bl_32 br_32 wl_120 vdd gnd cell_6t
Xbit_r121_c32 bl_32 br_32 wl_121 vdd gnd cell_6t
Xbit_r122_c32 bl_32 br_32 wl_122 vdd gnd cell_6t
Xbit_r123_c32 bl_32 br_32 wl_123 vdd gnd cell_6t
Xbit_r124_c32 bl_32 br_32 wl_124 vdd gnd cell_6t
Xbit_r125_c32 bl_32 br_32 wl_125 vdd gnd cell_6t
Xbit_r126_c32 bl_32 br_32 wl_126 vdd gnd cell_6t
Xbit_r127_c32 bl_32 br_32 wl_127 vdd gnd cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd cell_6t
Xbit_r1_c33 bl_33 br_33 wl_1 vdd gnd cell_6t
Xbit_r2_c33 bl_33 br_33 wl_2 vdd gnd cell_6t
Xbit_r3_c33 bl_33 br_33 wl_3 vdd gnd cell_6t
Xbit_r4_c33 bl_33 br_33 wl_4 vdd gnd cell_6t
Xbit_r5_c33 bl_33 br_33 wl_5 vdd gnd cell_6t
Xbit_r6_c33 bl_33 br_33 wl_6 vdd gnd cell_6t
Xbit_r7_c33 bl_33 br_33 wl_7 vdd gnd cell_6t
Xbit_r8_c33 bl_33 br_33 wl_8 vdd gnd cell_6t
Xbit_r9_c33 bl_33 br_33 wl_9 vdd gnd cell_6t
Xbit_r10_c33 bl_33 br_33 wl_10 vdd gnd cell_6t
Xbit_r11_c33 bl_33 br_33 wl_11 vdd gnd cell_6t
Xbit_r12_c33 bl_33 br_33 wl_12 vdd gnd cell_6t
Xbit_r13_c33 bl_33 br_33 wl_13 vdd gnd cell_6t
Xbit_r14_c33 bl_33 br_33 wl_14 vdd gnd cell_6t
Xbit_r15_c33 bl_33 br_33 wl_15 vdd gnd cell_6t
Xbit_r16_c33 bl_33 br_33 wl_16 vdd gnd cell_6t
Xbit_r17_c33 bl_33 br_33 wl_17 vdd gnd cell_6t
Xbit_r18_c33 bl_33 br_33 wl_18 vdd gnd cell_6t
Xbit_r19_c33 bl_33 br_33 wl_19 vdd gnd cell_6t
Xbit_r20_c33 bl_33 br_33 wl_20 vdd gnd cell_6t
Xbit_r21_c33 bl_33 br_33 wl_21 vdd gnd cell_6t
Xbit_r22_c33 bl_33 br_33 wl_22 vdd gnd cell_6t
Xbit_r23_c33 bl_33 br_33 wl_23 vdd gnd cell_6t
Xbit_r24_c33 bl_33 br_33 wl_24 vdd gnd cell_6t
Xbit_r25_c33 bl_33 br_33 wl_25 vdd gnd cell_6t
Xbit_r26_c33 bl_33 br_33 wl_26 vdd gnd cell_6t
Xbit_r27_c33 bl_33 br_33 wl_27 vdd gnd cell_6t
Xbit_r28_c33 bl_33 br_33 wl_28 vdd gnd cell_6t
Xbit_r29_c33 bl_33 br_33 wl_29 vdd gnd cell_6t
Xbit_r30_c33 bl_33 br_33 wl_30 vdd gnd cell_6t
Xbit_r31_c33 bl_33 br_33 wl_31 vdd gnd cell_6t
Xbit_r32_c33 bl_33 br_33 wl_32 vdd gnd cell_6t
Xbit_r33_c33 bl_33 br_33 wl_33 vdd gnd cell_6t
Xbit_r34_c33 bl_33 br_33 wl_34 vdd gnd cell_6t
Xbit_r35_c33 bl_33 br_33 wl_35 vdd gnd cell_6t
Xbit_r36_c33 bl_33 br_33 wl_36 vdd gnd cell_6t
Xbit_r37_c33 bl_33 br_33 wl_37 vdd gnd cell_6t
Xbit_r38_c33 bl_33 br_33 wl_38 vdd gnd cell_6t
Xbit_r39_c33 bl_33 br_33 wl_39 vdd gnd cell_6t
Xbit_r40_c33 bl_33 br_33 wl_40 vdd gnd cell_6t
Xbit_r41_c33 bl_33 br_33 wl_41 vdd gnd cell_6t
Xbit_r42_c33 bl_33 br_33 wl_42 vdd gnd cell_6t
Xbit_r43_c33 bl_33 br_33 wl_43 vdd gnd cell_6t
Xbit_r44_c33 bl_33 br_33 wl_44 vdd gnd cell_6t
Xbit_r45_c33 bl_33 br_33 wl_45 vdd gnd cell_6t
Xbit_r46_c33 bl_33 br_33 wl_46 vdd gnd cell_6t
Xbit_r47_c33 bl_33 br_33 wl_47 vdd gnd cell_6t
Xbit_r48_c33 bl_33 br_33 wl_48 vdd gnd cell_6t
Xbit_r49_c33 bl_33 br_33 wl_49 vdd gnd cell_6t
Xbit_r50_c33 bl_33 br_33 wl_50 vdd gnd cell_6t
Xbit_r51_c33 bl_33 br_33 wl_51 vdd gnd cell_6t
Xbit_r52_c33 bl_33 br_33 wl_52 vdd gnd cell_6t
Xbit_r53_c33 bl_33 br_33 wl_53 vdd gnd cell_6t
Xbit_r54_c33 bl_33 br_33 wl_54 vdd gnd cell_6t
Xbit_r55_c33 bl_33 br_33 wl_55 vdd gnd cell_6t
Xbit_r56_c33 bl_33 br_33 wl_56 vdd gnd cell_6t
Xbit_r57_c33 bl_33 br_33 wl_57 vdd gnd cell_6t
Xbit_r58_c33 bl_33 br_33 wl_58 vdd gnd cell_6t
Xbit_r59_c33 bl_33 br_33 wl_59 vdd gnd cell_6t
Xbit_r60_c33 bl_33 br_33 wl_60 vdd gnd cell_6t
Xbit_r61_c33 bl_33 br_33 wl_61 vdd gnd cell_6t
Xbit_r62_c33 bl_33 br_33 wl_62 vdd gnd cell_6t
Xbit_r63_c33 bl_33 br_33 wl_63 vdd gnd cell_6t
Xbit_r64_c33 bl_33 br_33 wl_64 vdd gnd cell_6t
Xbit_r65_c33 bl_33 br_33 wl_65 vdd gnd cell_6t
Xbit_r66_c33 bl_33 br_33 wl_66 vdd gnd cell_6t
Xbit_r67_c33 bl_33 br_33 wl_67 vdd gnd cell_6t
Xbit_r68_c33 bl_33 br_33 wl_68 vdd gnd cell_6t
Xbit_r69_c33 bl_33 br_33 wl_69 vdd gnd cell_6t
Xbit_r70_c33 bl_33 br_33 wl_70 vdd gnd cell_6t
Xbit_r71_c33 bl_33 br_33 wl_71 vdd gnd cell_6t
Xbit_r72_c33 bl_33 br_33 wl_72 vdd gnd cell_6t
Xbit_r73_c33 bl_33 br_33 wl_73 vdd gnd cell_6t
Xbit_r74_c33 bl_33 br_33 wl_74 vdd gnd cell_6t
Xbit_r75_c33 bl_33 br_33 wl_75 vdd gnd cell_6t
Xbit_r76_c33 bl_33 br_33 wl_76 vdd gnd cell_6t
Xbit_r77_c33 bl_33 br_33 wl_77 vdd gnd cell_6t
Xbit_r78_c33 bl_33 br_33 wl_78 vdd gnd cell_6t
Xbit_r79_c33 bl_33 br_33 wl_79 vdd gnd cell_6t
Xbit_r80_c33 bl_33 br_33 wl_80 vdd gnd cell_6t
Xbit_r81_c33 bl_33 br_33 wl_81 vdd gnd cell_6t
Xbit_r82_c33 bl_33 br_33 wl_82 vdd gnd cell_6t
Xbit_r83_c33 bl_33 br_33 wl_83 vdd gnd cell_6t
Xbit_r84_c33 bl_33 br_33 wl_84 vdd gnd cell_6t
Xbit_r85_c33 bl_33 br_33 wl_85 vdd gnd cell_6t
Xbit_r86_c33 bl_33 br_33 wl_86 vdd gnd cell_6t
Xbit_r87_c33 bl_33 br_33 wl_87 vdd gnd cell_6t
Xbit_r88_c33 bl_33 br_33 wl_88 vdd gnd cell_6t
Xbit_r89_c33 bl_33 br_33 wl_89 vdd gnd cell_6t
Xbit_r90_c33 bl_33 br_33 wl_90 vdd gnd cell_6t
Xbit_r91_c33 bl_33 br_33 wl_91 vdd gnd cell_6t
Xbit_r92_c33 bl_33 br_33 wl_92 vdd gnd cell_6t
Xbit_r93_c33 bl_33 br_33 wl_93 vdd gnd cell_6t
Xbit_r94_c33 bl_33 br_33 wl_94 vdd gnd cell_6t
Xbit_r95_c33 bl_33 br_33 wl_95 vdd gnd cell_6t
Xbit_r96_c33 bl_33 br_33 wl_96 vdd gnd cell_6t
Xbit_r97_c33 bl_33 br_33 wl_97 vdd gnd cell_6t
Xbit_r98_c33 bl_33 br_33 wl_98 vdd gnd cell_6t
Xbit_r99_c33 bl_33 br_33 wl_99 vdd gnd cell_6t
Xbit_r100_c33 bl_33 br_33 wl_100 vdd gnd cell_6t
Xbit_r101_c33 bl_33 br_33 wl_101 vdd gnd cell_6t
Xbit_r102_c33 bl_33 br_33 wl_102 vdd gnd cell_6t
Xbit_r103_c33 bl_33 br_33 wl_103 vdd gnd cell_6t
Xbit_r104_c33 bl_33 br_33 wl_104 vdd gnd cell_6t
Xbit_r105_c33 bl_33 br_33 wl_105 vdd gnd cell_6t
Xbit_r106_c33 bl_33 br_33 wl_106 vdd gnd cell_6t
Xbit_r107_c33 bl_33 br_33 wl_107 vdd gnd cell_6t
Xbit_r108_c33 bl_33 br_33 wl_108 vdd gnd cell_6t
Xbit_r109_c33 bl_33 br_33 wl_109 vdd gnd cell_6t
Xbit_r110_c33 bl_33 br_33 wl_110 vdd gnd cell_6t
Xbit_r111_c33 bl_33 br_33 wl_111 vdd gnd cell_6t
Xbit_r112_c33 bl_33 br_33 wl_112 vdd gnd cell_6t
Xbit_r113_c33 bl_33 br_33 wl_113 vdd gnd cell_6t
Xbit_r114_c33 bl_33 br_33 wl_114 vdd gnd cell_6t
Xbit_r115_c33 bl_33 br_33 wl_115 vdd gnd cell_6t
Xbit_r116_c33 bl_33 br_33 wl_116 vdd gnd cell_6t
Xbit_r117_c33 bl_33 br_33 wl_117 vdd gnd cell_6t
Xbit_r118_c33 bl_33 br_33 wl_118 vdd gnd cell_6t
Xbit_r119_c33 bl_33 br_33 wl_119 vdd gnd cell_6t
Xbit_r120_c33 bl_33 br_33 wl_120 vdd gnd cell_6t
Xbit_r121_c33 bl_33 br_33 wl_121 vdd gnd cell_6t
Xbit_r122_c33 bl_33 br_33 wl_122 vdd gnd cell_6t
Xbit_r123_c33 bl_33 br_33 wl_123 vdd gnd cell_6t
Xbit_r124_c33 bl_33 br_33 wl_124 vdd gnd cell_6t
Xbit_r125_c33 bl_33 br_33 wl_125 vdd gnd cell_6t
Xbit_r126_c33 bl_33 br_33 wl_126 vdd gnd cell_6t
Xbit_r127_c33 bl_33 br_33 wl_127 vdd gnd cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd cell_6t
Xbit_r1_c34 bl_34 br_34 wl_1 vdd gnd cell_6t
Xbit_r2_c34 bl_34 br_34 wl_2 vdd gnd cell_6t
Xbit_r3_c34 bl_34 br_34 wl_3 vdd gnd cell_6t
Xbit_r4_c34 bl_34 br_34 wl_4 vdd gnd cell_6t
Xbit_r5_c34 bl_34 br_34 wl_5 vdd gnd cell_6t
Xbit_r6_c34 bl_34 br_34 wl_6 vdd gnd cell_6t
Xbit_r7_c34 bl_34 br_34 wl_7 vdd gnd cell_6t
Xbit_r8_c34 bl_34 br_34 wl_8 vdd gnd cell_6t
Xbit_r9_c34 bl_34 br_34 wl_9 vdd gnd cell_6t
Xbit_r10_c34 bl_34 br_34 wl_10 vdd gnd cell_6t
Xbit_r11_c34 bl_34 br_34 wl_11 vdd gnd cell_6t
Xbit_r12_c34 bl_34 br_34 wl_12 vdd gnd cell_6t
Xbit_r13_c34 bl_34 br_34 wl_13 vdd gnd cell_6t
Xbit_r14_c34 bl_34 br_34 wl_14 vdd gnd cell_6t
Xbit_r15_c34 bl_34 br_34 wl_15 vdd gnd cell_6t
Xbit_r16_c34 bl_34 br_34 wl_16 vdd gnd cell_6t
Xbit_r17_c34 bl_34 br_34 wl_17 vdd gnd cell_6t
Xbit_r18_c34 bl_34 br_34 wl_18 vdd gnd cell_6t
Xbit_r19_c34 bl_34 br_34 wl_19 vdd gnd cell_6t
Xbit_r20_c34 bl_34 br_34 wl_20 vdd gnd cell_6t
Xbit_r21_c34 bl_34 br_34 wl_21 vdd gnd cell_6t
Xbit_r22_c34 bl_34 br_34 wl_22 vdd gnd cell_6t
Xbit_r23_c34 bl_34 br_34 wl_23 vdd gnd cell_6t
Xbit_r24_c34 bl_34 br_34 wl_24 vdd gnd cell_6t
Xbit_r25_c34 bl_34 br_34 wl_25 vdd gnd cell_6t
Xbit_r26_c34 bl_34 br_34 wl_26 vdd gnd cell_6t
Xbit_r27_c34 bl_34 br_34 wl_27 vdd gnd cell_6t
Xbit_r28_c34 bl_34 br_34 wl_28 vdd gnd cell_6t
Xbit_r29_c34 bl_34 br_34 wl_29 vdd gnd cell_6t
Xbit_r30_c34 bl_34 br_34 wl_30 vdd gnd cell_6t
Xbit_r31_c34 bl_34 br_34 wl_31 vdd gnd cell_6t
Xbit_r32_c34 bl_34 br_34 wl_32 vdd gnd cell_6t
Xbit_r33_c34 bl_34 br_34 wl_33 vdd gnd cell_6t
Xbit_r34_c34 bl_34 br_34 wl_34 vdd gnd cell_6t
Xbit_r35_c34 bl_34 br_34 wl_35 vdd gnd cell_6t
Xbit_r36_c34 bl_34 br_34 wl_36 vdd gnd cell_6t
Xbit_r37_c34 bl_34 br_34 wl_37 vdd gnd cell_6t
Xbit_r38_c34 bl_34 br_34 wl_38 vdd gnd cell_6t
Xbit_r39_c34 bl_34 br_34 wl_39 vdd gnd cell_6t
Xbit_r40_c34 bl_34 br_34 wl_40 vdd gnd cell_6t
Xbit_r41_c34 bl_34 br_34 wl_41 vdd gnd cell_6t
Xbit_r42_c34 bl_34 br_34 wl_42 vdd gnd cell_6t
Xbit_r43_c34 bl_34 br_34 wl_43 vdd gnd cell_6t
Xbit_r44_c34 bl_34 br_34 wl_44 vdd gnd cell_6t
Xbit_r45_c34 bl_34 br_34 wl_45 vdd gnd cell_6t
Xbit_r46_c34 bl_34 br_34 wl_46 vdd gnd cell_6t
Xbit_r47_c34 bl_34 br_34 wl_47 vdd gnd cell_6t
Xbit_r48_c34 bl_34 br_34 wl_48 vdd gnd cell_6t
Xbit_r49_c34 bl_34 br_34 wl_49 vdd gnd cell_6t
Xbit_r50_c34 bl_34 br_34 wl_50 vdd gnd cell_6t
Xbit_r51_c34 bl_34 br_34 wl_51 vdd gnd cell_6t
Xbit_r52_c34 bl_34 br_34 wl_52 vdd gnd cell_6t
Xbit_r53_c34 bl_34 br_34 wl_53 vdd gnd cell_6t
Xbit_r54_c34 bl_34 br_34 wl_54 vdd gnd cell_6t
Xbit_r55_c34 bl_34 br_34 wl_55 vdd gnd cell_6t
Xbit_r56_c34 bl_34 br_34 wl_56 vdd gnd cell_6t
Xbit_r57_c34 bl_34 br_34 wl_57 vdd gnd cell_6t
Xbit_r58_c34 bl_34 br_34 wl_58 vdd gnd cell_6t
Xbit_r59_c34 bl_34 br_34 wl_59 vdd gnd cell_6t
Xbit_r60_c34 bl_34 br_34 wl_60 vdd gnd cell_6t
Xbit_r61_c34 bl_34 br_34 wl_61 vdd gnd cell_6t
Xbit_r62_c34 bl_34 br_34 wl_62 vdd gnd cell_6t
Xbit_r63_c34 bl_34 br_34 wl_63 vdd gnd cell_6t
Xbit_r64_c34 bl_34 br_34 wl_64 vdd gnd cell_6t
Xbit_r65_c34 bl_34 br_34 wl_65 vdd gnd cell_6t
Xbit_r66_c34 bl_34 br_34 wl_66 vdd gnd cell_6t
Xbit_r67_c34 bl_34 br_34 wl_67 vdd gnd cell_6t
Xbit_r68_c34 bl_34 br_34 wl_68 vdd gnd cell_6t
Xbit_r69_c34 bl_34 br_34 wl_69 vdd gnd cell_6t
Xbit_r70_c34 bl_34 br_34 wl_70 vdd gnd cell_6t
Xbit_r71_c34 bl_34 br_34 wl_71 vdd gnd cell_6t
Xbit_r72_c34 bl_34 br_34 wl_72 vdd gnd cell_6t
Xbit_r73_c34 bl_34 br_34 wl_73 vdd gnd cell_6t
Xbit_r74_c34 bl_34 br_34 wl_74 vdd gnd cell_6t
Xbit_r75_c34 bl_34 br_34 wl_75 vdd gnd cell_6t
Xbit_r76_c34 bl_34 br_34 wl_76 vdd gnd cell_6t
Xbit_r77_c34 bl_34 br_34 wl_77 vdd gnd cell_6t
Xbit_r78_c34 bl_34 br_34 wl_78 vdd gnd cell_6t
Xbit_r79_c34 bl_34 br_34 wl_79 vdd gnd cell_6t
Xbit_r80_c34 bl_34 br_34 wl_80 vdd gnd cell_6t
Xbit_r81_c34 bl_34 br_34 wl_81 vdd gnd cell_6t
Xbit_r82_c34 bl_34 br_34 wl_82 vdd gnd cell_6t
Xbit_r83_c34 bl_34 br_34 wl_83 vdd gnd cell_6t
Xbit_r84_c34 bl_34 br_34 wl_84 vdd gnd cell_6t
Xbit_r85_c34 bl_34 br_34 wl_85 vdd gnd cell_6t
Xbit_r86_c34 bl_34 br_34 wl_86 vdd gnd cell_6t
Xbit_r87_c34 bl_34 br_34 wl_87 vdd gnd cell_6t
Xbit_r88_c34 bl_34 br_34 wl_88 vdd gnd cell_6t
Xbit_r89_c34 bl_34 br_34 wl_89 vdd gnd cell_6t
Xbit_r90_c34 bl_34 br_34 wl_90 vdd gnd cell_6t
Xbit_r91_c34 bl_34 br_34 wl_91 vdd gnd cell_6t
Xbit_r92_c34 bl_34 br_34 wl_92 vdd gnd cell_6t
Xbit_r93_c34 bl_34 br_34 wl_93 vdd gnd cell_6t
Xbit_r94_c34 bl_34 br_34 wl_94 vdd gnd cell_6t
Xbit_r95_c34 bl_34 br_34 wl_95 vdd gnd cell_6t
Xbit_r96_c34 bl_34 br_34 wl_96 vdd gnd cell_6t
Xbit_r97_c34 bl_34 br_34 wl_97 vdd gnd cell_6t
Xbit_r98_c34 bl_34 br_34 wl_98 vdd gnd cell_6t
Xbit_r99_c34 bl_34 br_34 wl_99 vdd gnd cell_6t
Xbit_r100_c34 bl_34 br_34 wl_100 vdd gnd cell_6t
Xbit_r101_c34 bl_34 br_34 wl_101 vdd gnd cell_6t
Xbit_r102_c34 bl_34 br_34 wl_102 vdd gnd cell_6t
Xbit_r103_c34 bl_34 br_34 wl_103 vdd gnd cell_6t
Xbit_r104_c34 bl_34 br_34 wl_104 vdd gnd cell_6t
Xbit_r105_c34 bl_34 br_34 wl_105 vdd gnd cell_6t
Xbit_r106_c34 bl_34 br_34 wl_106 vdd gnd cell_6t
Xbit_r107_c34 bl_34 br_34 wl_107 vdd gnd cell_6t
Xbit_r108_c34 bl_34 br_34 wl_108 vdd gnd cell_6t
Xbit_r109_c34 bl_34 br_34 wl_109 vdd gnd cell_6t
Xbit_r110_c34 bl_34 br_34 wl_110 vdd gnd cell_6t
Xbit_r111_c34 bl_34 br_34 wl_111 vdd gnd cell_6t
Xbit_r112_c34 bl_34 br_34 wl_112 vdd gnd cell_6t
Xbit_r113_c34 bl_34 br_34 wl_113 vdd gnd cell_6t
Xbit_r114_c34 bl_34 br_34 wl_114 vdd gnd cell_6t
Xbit_r115_c34 bl_34 br_34 wl_115 vdd gnd cell_6t
Xbit_r116_c34 bl_34 br_34 wl_116 vdd gnd cell_6t
Xbit_r117_c34 bl_34 br_34 wl_117 vdd gnd cell_6t
Xbit_r118_c34 bl_34 br_34 wl_118 vdd gnd cell_6t
Xbit_r119_c34 bl_34 br_34 wl_119 vdd gnd cell_6t
Xbit_r120_c34 bl_34 br_34 wl_120 vdd gnd cell_6t
Xbit_r121_c34 bl_34 br_34 wl_121 vdd gnd cell_6t
Xbit_r122_c34 bl_34 br_34 wl_122 vdd gnd cell_6t
Xbit_r123_c34 bl_34 br_34 wl_123 vdd gnd cell_6t
Xbit_r124_c34 bl_34 br_34 wl_124 vdd gnd cell_6t
Xbit_r125_c34 bl_34 br_34 wl_125 vdd gnd cell_6t
Xbit_r126_c34 bl_34 br_34 wl_126 vdd gnd cell_6t
Xbit_r127_c34 bl_34 br_34 wl_127 vdd gnd cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd cell_6t
Xbit_r1_c35 bl_35 br_35 wl_1 vdd gnd cell_6t
Xbit_r2_c35 bl_35 br_35 wl_2 vdd gnd cell_6t
Xbit_r3_c35 bl_35 br_35 wl_3 vdd gnd cell_6t
Xbit_r4_c35 bl_35 br_35 wl_4 vdd gnd cell_6t
Xbit_r5_c35 bl_35 br_35 wl_5 vdd gnd cell_6t
Xbit_r6_c35 bl_35 br_35 wl_6 vdd gnd cell_6t
Xbit_r7_c35 bl_35 br_35 wl_7 vdd gnd cell_6t
Xbit_r8_c35 bl_35 br_35 wl_8 vdd gnd cell_6t
Xbit_r9_c35 bl_35 br_35 wl_9 vdd gnd cell_6t
Xbit_r10_c35 bl_35 br_35 wl_10 vdd gnd cell_6t
Xbit_r11_c35 bl_35 br_35 wl_11 vdd gnd cell_6t
Xbit_r12_c35 bl_35 br_35 wl_12 vdd gnd cell_6t
Xbit_r13_c35 bl_35 br_35 wl_13 vdd gnd cell_6t
Xbit_r14_c35 bl_35 br_35 wl_14 vdd gnd cell_6t
Xbit_r15_c35 bl_35 br_35 wl_15 vdd gnd cell_6t
Xbit_r16_c35 bl_35 br_35 wl_16 vdd gnd cell_6t
Xbit_r17_c35 bl_35 br_35 wl_17 vdd gnd cell_6t
Xbit_r18_c35 bl_35 br_35 wl_18 vdd gnd cell_6t
Xbit_r19_c35 bl_35 br_35 wl_19 vdd gnd cell_6t
Xbit_r20_c35 bl_35 br_35 wl_20 vdd gnd cell_6t
Xbit_r21_c35 bl_35 br_35 wl_21 vdd gnd cell_6t
Xbit_r22_c35 bl_35 br_35 wl_22 vdd gnd cell_6t
Xbit_r23_c35 bl_35 br_35 wl_23 vdd gnd cell_6t
Xbit_r24_c35 bl_35 br_35 wl_24 vdd gnd cell_6t
Xbit_r25_c35 bl_35 br_35 wl_25 vdd gnd cell_6t
Xbit_r26_c35 bl_35 br_35 wl_26 vdd gnd cell_6t
Xbit_r27_c35 bl_35 br_35 wl_27 vdd gnd cell_6t
Xbit_r28_c35 bl_35 br_35 wl_28 vdd gnd cell_6t
Xbit_r29_c35 bl_35 br_35 wl_29 vdd gnd cell_6t
Xbit_r30_c35 bl_35 br_35 wl_30 vdd gnd cell_6t
Xbit_r31_c35 bl_35 br_35 wl_31 vdd gnd cell_6t
Xbit_r32_c35 bl_35 br_35 wl_32 vdd gnd cell_6t
Xbit_r33_c35 bl_35 br_35 wl_33 vdd gnd cell_6t
Xbit_r34_c35 bl_35 br_35 wl_34 vdd gnd cell_6t
Xbit_r35_c35 bl_35 br_35 wl_35 vdd gnd cell_6t
Xbit_r36_c35 bl_35 br_35 wl_36 vdd gnd cell_6t
Xbit_r37_c35 bl_35 br_35 wl_37 vdd gnd cell_6t
Xbit_r38_c35 bl_35 br_35 wl_38 vdd gnd cell_6t
Xbit_r39_c35 bl_35 br_35 wl_39 vdd gnd cell_6t
Xbit_r40_c35 bl_35 br_35 wl_40 vdd gnd cell_6t
Xbit_r41_c35 bl_35 br_35 wl_41 vdd gnd cell_6t
Xbit_r42_c35 bl_35 br_35 wl_42 vdd gnd cell_6t
Xbit_r43_c35 bl_35 br_35 wl_43 vdd gnd cell_6t
Xbit_r44_c35 bl_35 br_35 wl_44 vdd gnd cell_6t
Xbit_r45_c35 bl_35 br_35 wl_45 vdd gnd cell_6t
Xbit_r46_c35 bl_35 br_35 wl_46 vdd gnd cell_6t
Xbit_r47_c35 bl_35 br_35 wl_47 vdd gnd cell_6t
Xbit_r48_c35 bl_35 br_35 wl_48 vdd gnd cell_6t
Xbit_r49_c35 bl_35 br_35 wl_49 vdd gnd cell_6t
Xbit_r50_c35 bl_35 br_35 wl_50 vdd gnd cell_6t
Xbit_r51_c35 bl_35 br_35 wl_51 vdd gnd cell_6t
Xbit_r52_c35 bl_35 br_35 wl_52 vdd gnd cell_6t
Xbit_r53_c35 bl_35 br_35 wl_53 vdd gnd cell_6t
Xbit_r54_c35 bl_35 br_35 wl_54 vdd gnd cell_6t
Xbit_r55_c35 bl_35 br_35 wl_55 vdd gnd cell_6t
Xbit_r56_c35 bl_35 br_35 wl_56 vdd gnd cell_6t
Xbit_r57_c35 bl_35 br_35 wl_57 vdd gnd cell_6t
Xbit_r58_c35 bl_35 br_35 wl_58 vdd gnd cell_6t
Xbit_r59_c35 bl_35 br_35 wl_59 vdd gnd cell_6t
Xbit_r60_c35 bl_35 br_35 wl_60 vdd gnd cell_6t
Xbit_r61_c35 bl_35 br_35 wl_61 vdd gnd cell_6t
Xbit_r62_c35 bl_35 br_35 wl_62 vdd gnd cell_6t
Xbit_r63_c35 bl_35 br_35 wl_63 vdd gnd cell_6t
Xbit_r64_c35 bl_35 br_35 wl_64 vdd gnd cell_6t
Xbit_r65_c35 bl_35 br_35 wl_65 vdd gnd cell_6t
Xbit_r66_c35 bl_35 br_35 wl_66 vdd gnd cell_6t
Xbit_r67_c35 bl_35 br_35 wl_67 vdd gnd cell_6t
Xbit_r68_c35 bl_35 br_35 wl_68 vdd gnd cell_6t
Xbit_r69_c35 bl_35 br_35 wl_69 vdd gnd cell_6t
Xbit_r70_c35 bl_35 br_35 wl_70 vdd gnd cell_6t
Xbit_r71_c35 bl_35 br_35 wl_71 vdd gnd cell_6t
Xbit_r72_c35 bl_35 br_35 wl_72 vdd gnd cell_6t
Xbit_r73_c35 bl_35 br_35 wl_73 vdd gnd cell_6t
Xbit_r74_c35 bl_35 br_35 wl_74 vdd gnd cell_6t
Xbit_r75_c35 bl_35 br_35 wl_75 vdd gnd cell_6t
Xbit_r76_c35 bl_35 br_35 wl_76 vdd gnd cell_6t
Xbit_r77_c35 bl_35 br_35 wl_77 vdd gnd cell_6t
Xbit_r78_c35 bl_35 br_35 wl_78 vdd gnd cell_6t
Xbit_r79_c35 bl_35 br_35 wl_79 vdd gnd cell_6t
Xbit_r80_c35 bl_35 br_35 wl_80 vdd gnd cell_6t
Xbit_r81_c35 bl_35 br_35 wl_81 vdd gnd cell_6t
Xbit_r82_c35 bl_35 br_35 wl_82 vdd gnd cell_6t
Xbit_r83_c35 bl_35 br_35 wl_83 vdd gnd cell_6t
Xbit_r84_c35 bl_35 br_35 wl_84 vdd gnd cell_6t
Xbit_r85_c35 bl_35 br_35 wl_85 vdd gnd cell_6t
Xbit_r86_c35 bl_35 br_35 wl_86 vdd gnd cell_6t
Xbit_r87_c35 bl_35 br_35 wl_87 vdd gnd cell_6t
Xbit_r88_c35 bl_35 br_35 wl_88 vdd gnd cell_6t
Xbit_r89_c35 bl_35 br_35 wl_89 vdd gnd cell_6t
Xbit_r90_c35 bl_35 br_35 wl_90 vdd gnd cell_6t
Xbit_r91_c35 bl_35 br_35 wl_91 vdd gnd cell_6t
Xbit_r92_c35 bl_35 br_35 wl_92 vdd gnd cell_6t
Xbit_r93_c35 bl_35 br_35 wl_93 vdd gnd cell_6t
Xbit_r94_c35 bl_35 br_35 wl_94 vdd gnd cell_6t
Xbit_r95_c35 bl_35 br_35 wl_95 vdd gnd cell_6t
Xbit_r96_c35 bl_35 br_35 wl_96 vdd gnd cell_6t
Xbit_r97_c35 bl_35 br_35 wl_97 vdd gnd cell_6t
Xbit_r98_c35 bl_35 br_35 wl_98 vdd gnd cell_6t
Xbit_r99_c35 bl_35 br_35 wl_99 vdd gnd cell_6t
Xbit_r100_c35 bl_35 br_35 wl_100 vdd gnd cell_6t
Xbit_r101_c35 bl_35 br_35 wl_101 vdd gnd cell_6t
Xbit_r102_c35 bl_35 br_35 wl_102 vdd gnd cell_6t
Xbit_r103_c35 bl_35 br_35 wl_103 vdd gnd cell_6t
Xbit_r104_c35 bl_35 br_35 wl_104 vdd gnd cell_6t
Xbit_r105_c35 bl_35 br_35 wl_105 vdd gnd cell_6t
Xbit_r106_c35 bl_35 br_35 wl_106 vdd gnd cell_6t
Xbit_r107_c35 bl_35 br_35 wl_107 vdd gnd cell_6t
Xbit_r108_c35 bl_35 br_35 wl_108 vdd gnd cell_6t
Xbit_r109_c35 bl_35 br_35 wl_109 vdd gnd cell_6t
Xbit_r110_c35 bl_35 br_35 wl_110 vdd gnd cell_6t
Xbit_r111_c35 bl_35 br_35 wl_111 vdd gnd cell_6t
Xbit_r112_c35 bl_35 br_35 wl_112 vdd gnd cell_6t
Xbit_r113_c35 bl_35 br_35 wl_113 vdd gnd cell_6t
Xbit_r114_c35 bl_35 br_35 wl_114 vdd gnd cell_6t
Xbit_r115_c35 bl_35 br_35 wl_115 vdd gnd cell_6t
Xbit_r116_c35 bl_35 br_35 wl_116 vdd gnd cell_6t
Xbit_r117_c35 bl_35 br_35 wl_117 vdd gnd cell_6t
Xbit_r118_c35 bl_35 br_35 wl_118 vdd gnd cell_6t
Xbit_r119_c35 bl_35 br_35 wl_119 vdd gnd cell_6t
Xbit_r120_c35 bl_35 br_35 wl_120 vdd gnd cell_6t
Xbit_r121_c35 bl_35 br_35 wl_121 vdd gnd cell_6t
Xbit_r122_c35 bl_35 br_35 wl_122 vdd gnd cell_6t
Xbit_r123_c35 bl_35 br_35 wl_123 vdd gnd cell_6t
Xbit_r124_c35 bl_35 br_35 wl_124 vdd gnd cell_6t
Xbit_r125_c35 bl_35 br_35 wl_125 vdd gnd cell_6t
Xbit_r126_c35 bl_35 br_35 wl_126 vdd gnd cell_6t
Xbit_r127_c35 bl_35 br_35 wl_127 vdd gnd cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd cell_6t
Xbit_r1_c36 bl_36 br_36 wl_1 vdd gnd cell_6t
Xbit_r2_c36 bl_36 br_36 wl_2 vdd gnd cell_6t
Xbit_r3_c36 bl_36 br_36 wl_3 vdd gnd cell_6t
Xbit_r4_c36 bl_36 br_36 wl_4 vdd gnd cell_6t
Xbit_r5_c36 bl_36 br_36 wl_5 vdd gnd cell_6t
Xbit_r6_c36 bl_36 br_36 wl_6 vdd gnd cell_6t
Xbit_r7_c36 bl_36 br_36 wl_7 vdd gnd cell_6t
Xbit_r8_c36 bl_36 br_36 wl_8 vdd gnd cell_6t
Xbit_r9_c36 bl_36 br_36 wl_9 vdd gnd cell_6t
Xbit_r10_c36 bl_36 br_36 wl_10 vdd gnd cell_6t
Xbit_r11_c36 bl_36 br_36 wl_11 vdd gnd cell_6t
Xbit_r12_c36 bl_36 br_36 wl_12 vdd gnd cell_6t
Xbit_r13_c36 bl_36 br_36 wl_13 vdd gnd cell_6t
Xbit_r14_c36 bl_36 br_36 wl_14 vdd gnd cell_6t
Xbit_r15_c36 bl_36 br_36 wl_15 vdd gnd cell_6t
Xbit_r16_c36 bl_36 br_36 wl_16 vdd gnd cell_6t
Xbit_r17_c36 bl_36 br_36 wl_17 vdd gnd cell_6t
Xbit_r18_c36 bl_36 br_36 wl_18 vdd gnd cell_6t
Xbit_r19_c36 bl_36 br_36 wl_19 vdd gnd cell_6t
Xbit_r20_c36 bl_36 br_36 wl_20 vdd gnd cell_6t
Xbit_r21_c36 bl_36 br_36 wl_21 vdd gnd cell_6t
Xbit_r22_c36 bl_36 br_36 wl_22 vdd gnd cell_6t
Xbit_r23_c36 bl_36 br_36 wl_23 vdd gnd cell_6t
Xbit_r24_c36 bl_36 br_36 wl_24 vdd gnd cell_6t
Xbit_r25_c36 bl_36 br_36 wl_25 vdd gnd cell_6t
Xbit_r26_c36 bl_36 br_36 wl_26 vdd gnd cell_6t
Xbit_r27_c36 bl_36 br_36 wl_27 vdd gnd cell_6t
Xbit_r28_c36 bl_36 br_36 wl_28 vdd gnd cell_6t
Xbit_r29_c36 bl_36 br_36 wl_29 vdd gnd cell_6t
Xbit_r30_c36 bl_36 br_36 wl_30 vdd gnd cell_6t
Xbit_r31_c36 bl_36 br_36 wl_31 vdd gnd cell_6t
Xbit_r32_c36 bl_36 br_36 wl_32 vdd gnd cell_6t
Xbit_r33_c36 bl_36 br_36 wl_33 vdd gnd cell_6t
Xbit_r34_c36 bl_36 br_36 wl_34 vdd gnd cell_6t
Xbit_r35_c36 bl_36 br_36 wl_35 vdd gnd cell_6t
Xbit_r36_c36 bl_36 br_36 wl_36 vdd gnd cell_6t
Xbit_r37_c36 bl_36 br_36 wl_37 vdd gnd cell_6t
Xbit_r38_c36 bl_36 br_36 wl_38 vdd gnd cell_6t
Xbit_r39_c36 bl_36 br_36 wl_39 vdd gnd cell_6t
Xbit_r40_c36 bl_36 br_36 wl_40 vdd gnd cell_6t
Xbit_r41_c36 bl_36 br_36 wl_41 vdd gnd cell_6t
Xbit_r42_c36 bl_36 br_36 wl_42 vdd gnd cell_6t
Xbit_r43_c36 bl_36 br_36 wl_43 vdd gnd cell_6t
Xbit_r44_c36 bl_36 br_36 wl_44 vdd gnd cell_6t
Xbit_r45_c36 bl_36 br_36 wl_45 vdd gnd cell_6t
Xbit_r46_c36 bl_36 br_36 wl_46 vdd gnd cell_6t
Xbit_r47_c36 bl_36 br_36 wl_47 vdd gnd cell_6t
Xbit_r48_c36 bl_36 br_36 wl_48 vdd gnd cell_6t
Xbit_r49_c36 bl_36 br_36 wl_49 vdd gnd cell_6t
Xbit_r50_c36 bl_36 br_36 wl_50 vdd gnd cell_6t
Xbit_r51_c36 bl_36 br_36 wl_51 vdd gnd cell_6t
Xbit_r52_c36 bl_36 br_36 wl_52 vdd gnd cell_6t
Xbit_r53_c36 bl_36 br_36 wl_53 vdd gnd cell_6t
Xbit_r54_c36 bl_36 br_36 wl_54 vdd gnd cell_6t
Xbit_r55_c36 bl_36 br_36 wl_55 vdd gnd cell_6t
Xbit_r56_c36 bl_36 br_36 wl_56 vdd gnd cell_6t
Xbit_r57_c36 bl_36 br_36 wl_57 vdd gnd cell_6t
Xbit_r58_c36 bl_36 br_36 wl_58 vdd gnd cell_6t
Xbit_r59_c36 bl_36 br_36 wl_59 vdd gnd cell_6t
Xbit_r60_c36 bl_36 br_36 wl_60 vdd gnd cell_6t
Xbit_r61_c36 bl_36 br_36 wl_61 vdd gnd cell_6t
Xbit_r62_c36 bl_36 br_36 wl_62 vdd gnd cell_6t
Xbit_r63_c36 bl_36 br_36 wl_63 vdd gnd cell_6t
Xbit_r64_c36 bl_36 br_36 wl_64 vdd gnd cell_6t
Xbit_r65_c36 bl_36 br_36 wl_65 vdd gnd cell_6t
Xbit_r66_c36 bl_36 br_36 wl_66 vdd gnd cell_6t
Xbit_r67_c36 bl_36 br_36 wl_67 vdd gnd cell_6t
Xbit_r68_c36 bl_36 br_36 wl_68 vdd gnd cell_6t
Xbit_r69_c36 bl_36 br_36 wl_69 vdd gnd cell_6t
Xbit_r70_c36 bl_36 br_36 wl_70 vdd gnd cell_6t
Xbit_r71_c36 bl_36 br_36 wl_71 vdd gnd cell_6t
Xbit_r72_c36 bl_36 br_36 wl_72 vdd gnd cell_6t
Xbit_r73_c36 bl_36 br_36 wl_73 vdd gnd cell_6t
Xbit_r74_c36 bl_36 br_36 wl_74 vdd gnd cell_6t
Xbit_r75_c36 bl_36 br_36 wl_75 vdd gnd cell_6t
Xbit_r76_c36 bl_36 br_36 wl_76 vdd gnd cell_6t
Xbit_r77_c36 bl_36 br_36 wl_77 vdd gnd cell_6t
Xbit_r78_c36 bl_36 br_36 wl_78 vdd gnd cell_6t
Xbit_r79_c36 bl_36 br_36 wl_79 vdd gnd cell_6t
Xbit_r80_c36 bl_36 br_36 wl_80 vdd gnd cell_6t
Xbit_r81_c36 bl_36 br_36 wl_81 vdd gnd cell_6t
Xbit_r82_c36 bl_36 br_36 wl_82 vdd gnd cell_6t
Xbit_r83_c36 bl_36 br_36 wl_83 vdd gnd cell_6t
Xbit_r84_c36 bl_36 br_36 wl_84 vdd gnd cell_6t
Xbit_r85_c36 bl_36 br_36 wl_85 vdd gnd cell_6t
Xbit_r86_c36 bl_36 br_36 wl_86 vdd gnd cell_6t
Xbit_r87_c36 bl_36 br_36 wl_87 vdd gnd cell_6t
Xbit_r88_c36 bl_36 br_36 wl_88 vdd gnd cell_6t
Xbit_r89_c36 bl_36 br_36 wl_89 vdd gnd cell_6t
Xbit_r90_c36 bl_36 br_36 wl_90 vdd gnd cell_6t
Xbit_r91_c36 bl_36 br_36 wl_91 vdd gnd cell_6t
Xbit_r92_c36 bl_36 br_36 wl_92 vdd gnd cell_6t
Xbit_r93_c36 bl_36 br_36 wl_93 vdd gnd cell_6t
Xbit_r94_c36 bl_36 br_36 wl_94 vdd gnd cell_6t
Xbit_r95_c36 bl_36 br_36 wl_95 vdd gnd cell_6t
Xbit_r96_c36 bl_36 br_36 wl_96 vdd gnd cell_6t
Xbit_r97_c36 bl_36 br_36 wl_97 vdd gnd cell_6t
Xbit_r98_c36 bl_36 br_36 wl_98 vdd gnd cell_6t
Xbit_r99_c36 bl_36 br_36 wl_99 vdd gnd cell_6t
Xbit_r100_c36 bl_36 br_36 wl_100 vdd gnd cell_6t
Xbit_r101_c36 bl_36 br_36 wl_101 vdd gnd cell_6t
Xbit_r102_c36 bl_36 br_36 wl_102 vdd gnd cell_6t
Xbit_r103_c36 bl_36 br_36 wl_103 vdd gnd cell_6t
Xbit_r104_c36 bl_36 br_36 wl_104 vdd gnd cell_6t
Xbit_r105_c36 bl_36 br_36 wl_105 vdd gnd cell_6t
Xbit_r106_c36 bl_36 br_36 wl_106 vdd gnd cell_6t
Xbit_r107_c36 bl_36 br_36 wl_107 vdd gnd cell_6t
Xbit_r108_c36 bl_36 br_36 wl_108 vdd gnd cell_6t
Xbit_r109_c36 bl_36 br_36 wl_109 vdd gnd cell_6t
Xbit_r110_c36 bl_36 br_36 wl_110 vdd gnd cell_6t
Xbit_r111_c36 bl_36 br_36 wl_111 vdd gnd cell_6t
Xbit_r112_c36 bl_36 br_36 wl_112 vdd gnd cell_6t
Xbit_r113_c36 bl_36 br_36 wl_113 vdd gnd cell_6t
Xbit_r114_c36 bl_36 br_36 wl_114 vdd gnd cell_6t
Xbit_r115_c36 bl_36 br_36 wl_115 vdd gnd cell_6t
Xbit_r116_c36 bl_36 br_36 wl_116 vdd gnd cell_6t
Xbit_r117_c36 bl_36 br_36 wl_117 vdd gnd cell_6t
Xbit_r118_c36 bl_36 br_36 wl_118 vdd gnd cell_6t
Xbit_r119_c36 bl_36 br_36 wl_119 vdd gnd cell_6t
Xbit_r120_c36 bl_36 br_36 wl_120 vdd gnd cell_6t
Xbit_r121_c36 bl_36 br_36 wl_121 vdd gnd cell_6t
Xbit_r122_c36 bl_36 br_36 wl_122 vdd gnd cell_6t
Xbit_r123_c36 bl_36 br_36 wl_123 vdd gnd cell_6t
Xbit_r124_c36 bl_36 br_36 wl_124 vdd gnd cell_6t
Xbit_r125_c36 bl_36 br_36 wl_125 vdd gnd cell_6t
Xbit_r126_c36 bl_36 br_36 wl_126 vdd gnd cell_6t
Xbit_r127_c36 bl_36 br_36 wl_127 vdd gnd cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd cell_6t
Xbit_r1_c37 bl_37 br_37 wl_1 vdd gnd cell_6t
Xbit_r2_c37 bl_37 br_37 wl_2 vdd gnd cell_6t
Xbit_r3_c37 bl_37 br_37 wl_3 vdd gnd cell_6t
Xbit_r4_c37 bl_37 br_37 wl_4 vdd gnd cell_6t
Xbit_r5_c37 bl_37 br_37 wl_5 vdd gnd cell_6t
Xbit_r6_c37 bl_37 br_37 wl_6 vdd gnd cell_6t
Xbit_r7_c37 bl_37 br_37 wl_7 vdd gnd cell_6t
Xbit_r8_c37 bl_37 br_37 wl_8 vdd gnd cell_6t
Xbit_r9_c37 bl_37 br_37 wl_9 vdd gnd cell_6t
Xbit_r10_c37 bl_37 br_37 wl_10 vdd gnd cell_6t
Xbit_r11_c37 bl_37 br_37 wl_11 vdd gnd cell_6t
Xbit_r12_c37 bl_37 br_37 wl_12 vdd gnd cell_6t
Xbit_r13_c37 bl_37 br_37 wl_13 vdd gnd cell_6t
Xbit_r14_c37 bl_37 br_37 wl_14 vdd gnd cell_6t
Xbit_r15_c37 bl_37 br_37 wl_15 vdd gnd cell_6t
Xbit_r16_c37 bl_37 br_37 wl_16 vdd gnd cell_6t
Xbit_r17_c37 bl_37 br_37 wl_17 vdd gnd cell_6t
Xbit_r18_c37 bl_37 br_37 wl_18 vdd gnd cell_6t
Xbit_r19_c37 bl_37 br_37 wl_19 vdd gnd cell_6t
Xbit_r20_c37 bl_37 br_37 wl_20 vdd gnd cell_6t
Xbit_r21_c37 bl_37 br_37 wl_21 vdd gnd cell_6t
Xbit_r22_c37 bl_37 br_37 wl_22 vdd gnd cell_6t
Xbit_r23_c37 bl_37 br_37 wl_23 vdd gnd cell_6t
Xbit_r24_c37 bl_37 br_37 wl_24 vdd gnd cell_6t
Xbit_r25_c37 bl_37 br_37 wl_25 vdd gnd cell_6t
Xbit_r26_c37 bl_37 br_37 wl_26 vdd gnd cell_6t
Xbit_r27_c37 bl_37 br_37 wl_27 vdd gnd cell_6t
Xbit_r28_c37 bl_37 br_37 wl_28 vdd gnd cell_6t
Xbit_r29_c37 bl_37 br_37 wl_29 vdd gnd cell_6t
Xbit_r30_c37 bl_37 br_37 wl_30 vdd gnd cell_6t
Xbit_r31_c37 bl_37 br_37 wl_31 vdd gnd cell_6t
Xbit_r32_c37 bl_37 br_37 wl_32 vdd gnd cell_6t
Xbit_r33_c37 bl_37 br_37 wl_33 vdd gnd cell_6t
Xbit_r34_c37 bl_37 br_37 wl_34 vdd gnd cell_6t
Xbit_r35_c37 bl_37 br_37 wl_35 vdd gnd cell_6t
Xbit_r36_c37 bl_37 br_37 wl_36 vdd gnd cell_6t
Xbit_r37_c37 bl_37 br_37 wl_37 vdd gnd cell_6t
Xbit_r38_c37 bl_37 br_37 wl_38 vdd gnd cell_6t
Xbit_r39_c37 bl_37 br_37 wl_39 vdd gnd cell_6t
Xbit_r40_c37 bl_37 br_37 wl_40 vdd gnd cell_6t
Xbit_r41_c37 bl_37 br_37 wl_41 vdd gnd cell_6t
Xbit_r42_c37 bl_37 br_37 wl_42 vdd gnd cell_6t
Xbit_r43_c37 bl_37 br_37 wl_43 vdd gnd cell_6t
Xbit_r44_c37 bl_37 br_37 wl_44 vdd gnd cell_6t
Xbit_r45_c37 bl_37 br_37 wl_45 vdd gnd cell_6t
Xbit_r46_c37 bl_37 br_37 wl_46 vdd gnd cell_6t
Xbit_r47_c37 bl_37 br_37 wl_47 vdd gnd cell_6t
Xbit_r48_c37 bl_37 br_37 wl_48 vdd gnd cell_6t
Xbit_r49_c37 bl_37 br_37 wl_49 vdd gnd cell_6t
Xbit_r50_c37 bl_37 br_37 wl_50 vdd gnd cell_6t
Xbit_r51_c37 bl_37 br_37 wl_51 vdd gnd cell_6t
Xbit_r52_c37 bl_37 br_37 wl_52 vdd gnd cell_6t
Xbit_r53_c37 bl_37 br_37 wl_53 vdd gnd cell_6t
Xbit_r54_c37 bl_37 br_37 wl_54 vdd gnd cell_6t
Xbit_r55_c37 bl_37 br_37 wl_55 vdd gnd cell_6t
Xbit_r56_c37 bl_37 br_37 wl_56 vdd gnd cell_6t
Xbit_r57_c37 bl_37 br_37 wl_57 vdd gnd cell_6t
Xbit_r58_c37 bl_37 br_37 wl_58 vdd gnd cell_6t
Xbit_r59_c37 bl_37 br_37 wl_59 vdd gnd cell_6t
Xbit_r60_c37 bl_37 br_37 wl_60 vdd gnd cell_6t
Xbit_r61_c37 bl_37 br_37 wl_61 vdd gnd cell_6t
Xbit_r62_c37 bl_37 br_37 wl_62 vdd gnd cell_6t
Xbit_r63_c37 bl_37 br_37 wl_63 vdd gnd cell_6t
Xbit_r64_c37 bl_37 br_37 wl_64 vdd gnd cell_6t
Xbit_r65_c37 bl_37 br_37 wl_65 vdd gnd cell_6t
Xbit_r66_c37 bl_37 br_37 wl_66 vdd gnd cell_6t
Xbit_r67_c37 bl_37 br_37 wl_67 vdd gnd cell_6t
Xbit_r68_c37 bl_37 br_37 wl_68 vdd gnd cell_6t
Xbit_r69_c37 bl_37 br_37 wl_69 vdd gnd cell_6t
Xbit_r70_c37 bl_37 br_37 wl_70 vdd gnd cell_6t
Xbit_r71_c37 bl_37 br_37 wl_71 vdd gnd cell_6t
Xbit_r72_c37 bl_37 br_37 wl_72 vdd gnd cell_6t
Xbit_r73_c37 bl_37 br_37 wl_73 vdd gnd cell_6t
Xbit_r74_c37 bl_37 br_37 wl_74 vdd gnd cell_6t
Xbit_r75_c37 bl_37 br_37 wl_75 vdd gnd cell_6t
Xbit_r76_c37 bl_37 br_37 wl_76 vdd gnd cell_6t
Xbit_r77_c37 bl_37 br_37 wl_77 vdd gnd cell_6t
Xbit_r78_c37 bl_37 br_37 wl_78 vdd gnd cell_6t
Xbit_r79_c37 bl_37 br_37 wl_79 vdd gnd cell_6t
Xbit_r80_c37 bl_37 br_37 wl_80 vdd gnd cell_6t
Xbit_r81_c37 bl_37 br_37 wl_81 vdd gnd cell_6t
Xbit_r82_c37 bl_37 br_37 wl_82 vdd gnd cell_6t
Xbit_r83_c37 bl_37 br_37 wl_83 vdd gnd cell_6t
Xbit_r84_c37 bl_37 br_37 wl_84 vdd gnd cell_6t
Xbit_r85_c37 bl_37 br_37 wl_85 vdd gnd cell_6t
Xbit_r86_c37 bl_37 br_37 wl_86 vdd gnd cell_6t
Xbit_r87_c37 bl_37 br_37 wl_87 vdd gnd cell_6t
Xbit_r88_c37 bl_37 br_37 wl_88 vdd gnd cell_6t
Xbit_r89_c37 bl_37 br_37 wl_89 vdd gnd cell_6t
Xbit_r90_c37 bl_37 br_37 wl_90 vdd gnd cell_6t
Xbit_r91_c37 bl_37 br_37 wl_91 vdd gnd cell_6t
Xbit_r92_c37 bl_37 br_37 wl_92 vdd gnd cell_6t
Xbit_r93_c37 bl_37 br_37 wl_93 vdd gnd cell_6t
Xbit_r94_c37 bl_37 br_37 wl_94 vdd gnd cell_6t
Xbit_r95_c37 bl_37 br_37 wl_95 vdd gnd cell_6t
Xbit_r96_c37 bl_37 br_37 wl_96 vdd gnd cell_6t
Xbit_r97_c37 bl_37 br_37 wl_97 vdd gnd cell_6t
Xbit_r98_c37 bl_37 br_37 wl_98 vdd gnd cell_6t
Xbit_r99_c37 bl_37 br_37 wl_99 vdd gnd cell_6t
Xbit_r100_c37 bl_37 br_37 wl_100 vdd gnd cell_6t
Xbit_r101_c37 bl_37 br_37 wl_101 vdd gnd cell_6t
Xbit_r102_c37 bl_37 br_37 wl_102 vdd gnd cell_6t
Xbit_r103_c37 bl_37 br_37 wl_103 vdd gnd cell_6t
Xbit_r104_c37 bl_37 br_37 wl_104 vdd gnd cell_6t
Xbit_r105_c37 bl_37 br_37 wl_105 vdd gnd cell_6t
Xbit_r106_c37 bl_37 br_37 wl_106 vdd gnd cell_6t
Xbit_r107_c37 bl_37 br_37 wl_107 vdd gnd cell_6t
Xbit_r108_c37 bl_37 br_37 wl_108 vdd gnd cell_6t
Xbit_r109_c37 bl_37 br_37 wl_109 vdd gnd cell_6t
Xbit_r110_c37 bl_37 br_37 wl_110 vdd gnd cell_6t
Xbit_r111_c37 bl_37 br_37 wl_111 vdd gnd cell_6t
Xbit_r112_c37 bl_37 br_37 wl_112 vdd gnd cell_6t
Xbit_r113_c37 bl_37 br_37 wl_113 vdd gnd cell_6t
Xbit_r114_c37 bl_37 br_37 wl_114 vdd gnd cell_6t
Xbit_r115_c37 bl_37 br_37 wl_115 vdd gnd cell_6t
Xbit_r116_c37 bl_37 br_37 wl_116 vdd gnd cell_6t
Xbit_r117_c37 bl_37 br_37 wl_117 vdd gnd cell_6t
Xbit_r118_c37 bl_37 br_37 wl_118 vdd gnd cell_6t
Xbit_r119_c37 bl_37 br_37 wl_119 vdd gnd cell_6t
Xbit_r120_c37 bl_37 br_37 wl_120 vdd gnd cell_6t
Xbit_r121_c37 bl_37 br_37 wl_121 vdd gnd cell_6t
Xbit_r122_c37 bl_37 br_37 wl_122 vdd gnd cell_6t
Xbit_r123_c37 bl_37 br_37 wl_123 vdd gnd cell_6t
Xbit_r124_c37 bl_37 br_37 wl_124 vdd gnd cell_6t
Xbit_r125_c37 bl_37 br_37 wl_125 vdd gnd cell_6t
Xbit_r126_c37 bl_37 br_37 wl_126 vdd gnd cell_6t
Xbit_r127_c37 bl_37 br_37 wl_127 vdd gnd cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd cell_6t
Xbit_r1_c38 bl_38 br_38 wl_1 vdd gnd cell_6t
Xbit_r2_c38 bl_38 br_38 wl_2 vdd gnd cell_6t
Xbit_r3_c38 bl_38 br_38 wl_3 vdd gnd cell_6t
Xbit_r4_c38 bl_38 br_38 wl_4 vdd gnd cell_6t
Xbit_r5_c38 bl_38 br_38 wl_5 vdd gnd cell_6t
Xbit_r6_c38 bl_38 br_38 wl_6 vdd gnd cell_6t
Xbit_r7_c38 bl_38 br_38 wl_7 vdd gnd cell_6t
Xbit_r8_c38 bl_38 br_38 wl_8 vdd gnd cell_6t
Xbit_r9_c38 bl_38 br_38 wl_9 vdd gnd cell_6t
Xbit_r10_c38 bl_38 br_38 wl_10 vdd gnd cell_6t
Xbit_r11_c38 bl_38 br_38 wl_11 vdd gnd cell_6t
Xbit_r12_c38 bl_38 br_38 wl_12 vdd gnd cell_6t
Xbit_r13_c38 bl_38 br_38 wl_13 vdd gnd cell_6t
Xbit_r14_c38 bl_38 br_38 wl_14 vdd gnd cell_6t
Xbit_r15_c38 bl_38 br_38 wl_15 vdd gnd cell_6t
Xbit_r16_c38 bl_38 br_38 wl_16 vdd gnd cell_6t
Xbit_r17_c38 bl_38 br_38 wl_17 vdd gnd cell_6t
Xbit_r18_c38 bl_38 br_38 wl_18 vdd gnd cell_6t
Xbit_r19_c38 bl_38 br_38 wl_19 vdd gnd cell_6t
Xbit_r20_c38 bl_38 br_38 wl_20 vdd gnd cell_6t
Xbit_r21_c38 bl_38 br_38 wl_21 vdd gnd cell_6t
Xbit_r22_c38 bl_38 br_38 wl_22 vdd gnd cell_6t
Xbit_r23_c38 bl_38 br_38 wl_23 vdd gnd cell_6t
Xbit_r24_c38 bl_38 br_38 wl_24 vdd gnd cell_6t
Xbit_r25_c38 bl_38 br_38 wl_25 vdd gnd cell_6t
Xbit_r26_c38 bl_38 br_38 wl_26 vdd gnd cell_6t
Xbit_r27_c38 bl_38 br_38 wl_27 vdd gnd cell_6t
Xbit_r28_c38 bl_38 br_38 wl_28 vdd gnd cell_6t
Xbit_r29_c38 bl_38 br_38 wl_29 vdd gnd cell_6t
Xbit_r30_c38 bl_38 br_38 wl_30 vdd gnd cell_6t
Xbit_r31_c38 bl_38 br_38 wl_31 vdd gnd cell_6t
Xbit_r32_c38 bl_38 br_38 wl_32 vdd gnd cell_6t
Xbit_r33_c38 bl_38 br_38 wl_33 vdd gnd cell_6t
Xbit_r34_c38 bl_38 br_38 wl_34 vdd gnd cell_6t
Xbit_r35_c38 bl_38 br_38 wl_35 vdd gnd cell_6t
Xbit_r36_c38 bl_38 br_38 wl_36 vdd gnd cell_6t
Xbit_r37_c38 bl_38 br_38 wl_37 vdd gnd cell_6t
Xbit_r38_c38 bl_38 br_38 wl_38 vdd gnd cell_6t
Xbit_r39_c38 bl_38 br_38 wl_39 vdd gnd cell_6t
Xbit_r40_c38 bl_38 br_38 wl_40 vdd gnd cell_6t
Xbit_r41_c38 bl_38 br_38 wl_41 vdd gnd cell_6t
Xbit_r42_c38 bl_38 br_38 wl_42 vdd gnd cell_6t
Xbit_r43_c38 bl_38 br_38 wl_43 vdd gnd cell_6t
Xbit_r44_c38 bl_38 br_38 wl_44 vdd gnd cell_6t
Xbit_r45_c38 bl_38 br_38 wl_45 vdd gnd cell_6t
Xbit_r46_c38 bl_38 br_38 wl_46 vdd gnd cell_6t
Xbit_r47_c38 bl_38 br_38 wl_47 vdd gnd cell_6t
Xbit_r48_c38 bl_38 br_38 wl_48 vdd gnd cell_6t
Xbit_r49_c38 bl_38 br_38 wl_49 vdd gnd cell_6t
Xbit_r50_c38 bl_38 br_38 wl_50 vdd gnd cell_6t
Xbit_r51_c38 bl_38 br_38 wl_51 vdd gnd cell_6t
Xbit_r52_c38 bl_38 br_38 wl_52 vdd gnd cell_6t
Xbit_r53_c38 bl_38 br_38 wl_53 vdd gnd cell_6t
Xbit_r54_c38 bl_38 br_38 wl_54 vdd gnd cell_6t
Xbit_r55_c38 bl_38 br_38 wl_55 vdd gnd cell_6t
Xbit_r56_c38 bl_38 br_38 wl_56 vdd gnd cell_6t
Xbit_r57_c38 bl_38 br_38 wl_57 vdd gnd cell_6t
Xbit_r58_c38 bl_38 br_38 wl_58 vdd gnd cell_6t
Xbit_r59_c38 bl_38 br_38 wl_59 vdd gnd cell_6t
Xbit_r60_c38 bl_38 br_38 wl_60 vdd gnd cell_6t
Xbit_r61_c38 bl_38 br_38 wl_61 vdd gnd cell_6t
Xbit_r62_c38 bl_38 br_38 wl_62 vdd gnd cell_6t
Xbit_r63_c38 bl_38 br_38 wl_63 vdd gnd cell_6t
Xbit_r64_c38 bl_38 br_38 wl_64 vdd gnd cell_6t
Xbit_r65_c38 bl_38 br_38 wl_65 vdd gnd cell_6t
Xbit_r66_c38 bl_38 br_38 wl_66 vdd gnd cell_6t
Xbit_r67_c38 bl_38 br_38 wl_67 vdd gnd cell_6t
Xbit_r68_c38 bl_38 br_38 wl_68 vdd gnd cell_6t
Xbit_r69_c38 bl_38 br_38 wl_69 vdd gnd cell_6t
Xbit_r70_c38 bl_38 br_38 wl_70 vdd gnd cell_6t
Xbit_r71_c38 bl_38 br_38 wl_71 vdd gnd cell_6t
Xbit_r72_c38 bl_38 br_38 wl_72 vdd gnd cell_6t
Xbit_r73_c38 bl_38 br_38 wl_73 vdd gnd cell_6t
Xbit_r74_c38 bl_38 br_38 wl_74 vdd gnd cell_6t
Xbit_r75_c38 bl_38 br_38 wl_75 vdd gnd cell_6t
Xbit_r76_c38 bl_38 br_38 wl_76 vdd gnd cell_6t
Xbit_r77_c38 bl_38 br_38 wl_77 vdd gnd cell_6t
Xbit_r78_c38 bl_38 br_38 wl_78 vdd gnd cell_6t
Xbit_r79_c38 bl_38 br_38 wl_79 vdd gnd cell_6t
Xbit_r80_c38 bl_38 br_38 wl_80 vdd gnd cell_6t
Xbit_r81_c38 bl_38 br_38 wl_81 vdd gnd cell_6t
Xbit_r82_c38 bl_38 br_38 wl_82 vdd gnd cell_6t
Xbit_r83_c38 bl_38 br_38 wl_83 vdd gnd cell_6t
Xbit_r84_c38 bl_38 br_38 wl_84 vdd gnd cell_6t
Xbit_r85_c38 bl_38 br_38 wl_85 vdd gnd cell_6t
Xbit_r86_c38 bl_38 br_38 wl_86 vdd gnd cell_6t
Xbit_r87_c38 bl_38 br_38 wl_87 vdd gnd cell_6t
Xbit_r88_c38 bl_38 br_38 wl_88 vdd gnd cell_6t
Xbit_r89_c38 bl_38 br_38 wl_89 vdd gnd cell_6t
Xbit_r90_c38 bl_38 br_38 wl_90 vdd gnd cell_6t
Xbit_r91_c38 bl_38 br_38 wl_91 vdd gnd cell_6t
Xbit_r92_c38 bl_38 br_38 wl_92 vdd gnd cell_6t
Xbit_r93_c38 bl_38 br_38 wl_93 vdd gnd cell_6t
Xbit_r94_c38 bl_38 br_38 wl_94 vdd gnd cell_6t
Xbit_r95_c38 bl_38 br_38 wl_95 vdd gnd cell_6t
Xbit_r96_c38 bl_38 br_38 wl_96 vdd gnd cell_6t
Xbit_r97_c38 bl_38 br_38 wl_97 vdd gnd cell_6t
Xbit_r98_c38 bl_38 br_38 wl_98 vdd gnd cell_6t
Xbit_r99_c38 bl_38 br_38 wl_99 vdd gnd cell_6t
Xbit_r100_c38 bl_38 br_38 wl_100 vdd gnd cell_6t
Xbit_r101_c38 bl_38 br_38 wl_101 vdd gnd cell_6t
Xbit_r102_c38 bl_38 br_38 wl_102 vdd gnd cell_6t
Xbit_r103_c38 bl_38 br_38 wl_103 vdd gnd cell_6t
Xbit_r104_c38 bl_38 br_38 wl_104 vdd gnd cell_6t
Xbit_r105_c38 bl_38 br_38 wl_105 vdd gnd cell_6t
Xbit_r106_c38 bl_38 br_38 wl_106 vdd gnd cell_6t
Xbit_r107_c38 bl_38 br_38 wl_107 vdd gnd cell_6t
Xbit_r108_c38 bl_38 br_38 wl_108 vdd gnd cell_6t
Xbit_r109_c38 bl_38 br_38 wl_109 vdd gnd cell_6t
Xbit_r110_c38 bl_38 br_38 wl_110 vdd gnd cell_6t
Xbit_r111_c38 bl_38 br_38 wl_111 vdd gnd cell_6t
Xbit_r112_c38 bl_38 br_38 wl_112 vdd gnd cell_6t
Xbit_r113_c38 bl_38 br_38 wl_113 vdd gnd cell_6t
Xbit_r114_c38 bl_38 br_38 wl_114 vdd gnd cell_6t
Xbit_r115_c38 bl_38 br_38 wl_115 vdd gnd cell_6t
Xbit_r116_c38 bl_38 br_38 wl_116 vdd gnd cell_6t
Xbit_r117_c38 bl_38 br_38 wl_117 vdd gnd cell_6t
Xbit_r118_c38 bl_38 br_38 wl_118 vdd gnd cell_6t
Xbit_r119_c38 bl_38 br_38 wl_119 vdd gnd cell_6t
Xbit_r120_c38 bl_38 br_38 wl_120 vdd gnd cell_6t
Xbit_r121_c38 bl_38 br_38 wl_121 vdd gnd cell_6t
Xbit_r122_c38 bl_38 br_38 wl_122 vdd gnd cell_6t
Xbit_r123_c38 bl_38 br_38 wl_123 vdd gnd cell_6t
Xbit_r124_c38 bl_38 br_38 wl_124 vdd gnd cell_6t
Xbit_r125_c38 bl_38 br_38 wl_125 vdd gnd cell_6t
Xbit_r126_c38 bl_38 br_38 wl_126 vdd gnd cell_6t
Xbit_r127_c38 bl_38 br_38 wl_127 vdd gnd cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd cell_6t
Xbit_r1_c39 bl_39 br_39 wl_1 vdd gnd cell_6t
Xbit_r2_c39 bl_39 br_39 wl_2 vdd gnd cell_6t
Xbit_r3_c39 bl_39 br_39 wl_3 vdd gnd cell_6t
Xbit_r4_c39 bl_39 br_39 wl_4 vdd gnd cell_6t
Xbit_r5_c39 bl_39 br_39 wl_5 vdd gnd cell_6t
Xbit_r6_c39 bl_39 br_39 wl_6 vdd gnd cell_6t
Xbit_r7_c39 bl_39 br_39 wl_7 vdd gnd cell_6t
Xbit_r8_c39 bl_39 br_39 wl_8 vdd gnd cell_6t
Xbit_r9_c39 bl_39 br_39 wl_9 vdd gnd cell_6t
Xbit_r10_c39 bl_39 br_39 wl_10 vdd gnd cell_6t
Xbit_r11_c39 bl_39 br_39 wl_11 vdd gnd cell_6t
Xbit_r12_c39 bl_39 br_39 wl_12 vdd gnd cell_6t
Xbit_r13_c39 bl_39 br_39 wl_13 vdd gnd cell_6t
Xbit_r14_c39 bl_39 br_39 wl_14 vdd gnd cell_6t
Xbit_r15_c39 bl_39 br_39 wl_15 vdd gnd cell_6t
Xbit_r16_c39 bl_39 br_39 wl_16 vdd gnd cell_6t
Xbit_r17_c39 bl_39 br_39 wl_17 vdd gnd cell_6t
Xbit_r18_c39 bl_39 br_39 wl_18 vdd gnd cell_6t
Xbit_r19_c39 bl_39 br_39 wl_19 vdd gnd cell_6t
Xbit_r20_c39 bl_39 br_39 wl_20 vdd gnd cell_6t
Xbit_r21_c39 bl_39 br_39 wl_21 vdd gnd cell_6t
Xbit_r22_c39 bl_39 br_39 wl_22 vdd gnd cell_6t
Xbit_r23_c39 bl_39 br_39 wl_23 vdd gnd cell_6t
Xbit_r24_c39 bl_39 br_39 wl_24 vdd gnd cell_6t
Xbit_r25_c39 bl_39 br_39 wl_25 vdd gnd cell_6t
Xbit_r26_c39 bl_39 br_39 wl_26 vdd gnd cell_6t
Xbit_r27_c39 bl_39 br_39 wl_27 vdd gnd cell_6t
Xbit_r28_c39 bl_39 br_39 wl_28 vdd gnd cell_6t
Xbit_r29_c39 bl_39 br_39 wl_29 vdd gnd cell_6t
Xbit_r30_c39 bl_39 br_39 wl_30 vdd gnd cell_6t
Xbit_r31_c39 bl_39 br_39 wl_31 vdd gnd cell_6t
Xbit_r32_c39 bl_39 br_39 wl_32 vdd gnd cell_6t
Xbit_r33_c39 bl_39 br_39 wl_33 vdd gnd cell_6t
Xbit_r34_c39 bl_39 br_39 wl_34 vdd gnd cell_6t
Xbit_r35_c39 bl_39 br_39 wl_35 vdd gnd cell_6t
Xbit_r36_c39 bl_39 br_39 wl_36 vdd gnd cell_6t
Xbit_r37_c39 bl_39 br_39 wl_37 vdd gnd cell_6t
Xbit_r38_c39 bl_39 br_39 wl_38 vdd gnd cell_6t
Xbit_r39_c39 bl_39 br_39 wl_39 vdd gnd cell_6t
Xbit_r40_c39 bl_39 br_39 wl_40 vdd gnd cell_6t
Xbit_r41_c39 bl_39 br_39 wl_41 vdd gnd cell_6t
Xbit_r42_c39 bl_39 br_39 wl_42 vdd gnd cell_6t
Xbit_r43_c39 bl_39 br_39 wl_43 vdd gnd cell_6t
Xbit_r44_c39 bl_39 br_39 wl_44 vdd gnd cell_6t
Xbit_r45_c39 bl_39 br_39 wl_45 vdd gnd cell_6t
Xbit_r46_c39 bl_39 br_39 wl_46 vdd gnd cell_6t
Xbit_r47_c39 bl_39 br_39 wl_47 vdd gnd cell_6t
Xbit_r48_c39 bl_39 br_39 wl_48 vdd gnd cell_6t
Xbit_r49_c39 bl_39 br_39 wl_49 vdd gnd cell_6t
Xbit_r50_c39 bl_39 br_39 wl_50 vdd gnd cell_6t
Xbit_r51_c39 bl_39 br_39 wl_51 vdd gnd cell_6t
Xbit_r52_c39 bl_39 br_39 wl_52 vdd gnd cell_6t
Xbit_r53_c39 bl_39 br_39 wl_53 vdd gnd cell_6t
Xbit_r54_c39 bl_39 br_39 wl_54 vdd gnd cell_6t
Xbit_r55_c39 bl_39 br_39 wl_55 vdd gnd cell_6t
Xbit_r56_c39 bl_39 br_39 wl_56 vdd gnd cell_6t
Xbit_r57_c39 bl_39 br_39 wl_57 vdd gnd cell_6t
Xbit_r58_c39 bl_39 br_39 wl_58 vdd gnd cell_6t
Xbit_r59_c39 bl_39 br_39 wl_59 vdd gnd cell_6t
Xbit_r60_c39 bl_39 br_39 wl_60 vdd gnd cell_6t
Xbit_r61_c39 bl_39 br_39 wl_61 vdd gnd cell_6t
Xbit_r62_c39 bl_39 br_39 wl_62 vdd gnd cell_6t
Xbit_r63_c39 bl_39 br_39 wl_63 vdd gnd cell_6t
Xbit_r64_c39 bl_39 br_39 wl_64 vdd gnd cell_6t
Xbit_r65_c39 bl_39 br_39 wl_65 vdd gnd cell_6t
Xbit_r66_c39 bl_39 br_39 wl_66 vdd gnd cell_6t
Xbit_r67_c39 bl_39 br_39 wl_67 vdd gnd cell_6t
Xbit_r68_c39 bl_39 br_39 wl_68 vdd gnd cell_6t
Xbit_r69_c39 bl_39 br_39 wl_69 vdd gnd cell_6t
Xbit_r70_c39 bl_39 br_39 wl_70 vdd gnd cell_6t
Xbit_r71_c39 bl_39 br_39 wl_71 vdd gnd cell_6t
Xbit_r72_c39 bl_39 br_39 wl_72 vdd gnd cell_6t
Xbit_r73_c39 bl_39 br_39 wl_73 vdd gnd cell_6t
Xbit_r74_c39 bl_39 br_39 wl_74 vdd gnd cell_6t
Xbit_r75_c39 bl_39 br_39 wl_75 vdd gnd cell_6t
Xbit_r76_c39 bl_39 br_39 wl_76 vdd gnd cell_6t
Xbit_r77_c39 bl_39 br_39 wl_77 vdd gnd cell_6t
Xbit_r78_c39 bl_39 br_39 wl_78 vdd gnd cell_6t
Xbit_r79_c39 bl_39 br_39 wl_79 vdd gnd cell_6t
Xbit_r80_c39 bl_39 br_39 wl_80 vdd gnd cell_6t
Xbit_r81_c39 bl_39 br_39 wl_81 vdd gnd cell_6t
Xbit_r82_c39 bl_39 br_39 wl_82 vdd gnd cell_6t
Xbit_r83_c39 bl_39 br_39 wl_83 vdd gnd cell_6t
Xbit_r84_c39 bl_39 br_39 wl_84 vdd gnd cell_6t
Xbit_r85_c39 bl_39 br_39 wl_85 vdd gnd cell_6t
Xbit_r86_c39 bl_39 br_39 wl_86 vdd gnd cell_6t
Xbit_r87_c39 bl_39 br_39 wl_87 vdd gnd cell_6t
Xbit_r88_c39 bl_39 br_39 wl_88 vdd gnd cell_6t
Xbit_r89_c39 bl_39 br_39 wl_89 vdd gnd cell_6t
Xbit_r90_c39 bl_39 br_39 wl_90 vdd gnd cell_6t
Xbit_r91_c39 bl_39 br_39 wl_91 vdd gnd cell_6t
Xbit_r92_c39 bl_39 br_39 wl_92 vdd gnd cell_6t
Xbit_r93_c39 bl_39 br_39 wl_93 vdd gnd cell_6t
Xbit_r94_c39 bl_39 br_39 wl_94 vdd gnd cell_6t
Xbit_r95_c39 bl_39 br_39 wl_95 vdd gnd cell_6t
Xbit_r96_c39 bl_39 br_39 wl_96 vdd gnd cell_6t
Xbit_r97_c39 bl_39 br_39 wl_97 vdd gnd cell_6t
Xbit_r98_c39 bl_39 br_39 wl_98 vdd gnd cell_6t
Xbit_r99_c39 bl_39 br_39 wl_99 vdd gnd cell_6t
Xbit_r100_c39 bl_39 br_39 wl_100 vdd gnd cell_6t
Xbit_r101_c39 bl_39 br_39 wl_101 vdd gnd cell_6t
Xbit_r102_c39 bl_39 br_39 wl_102 vdd gnd cell_6t
Xbit_r103_c39 bl_39 br_39 wl_103 vdd gnd cell_6t
Xbit_r104_c39 bl_39 br_39 wl_104 vdd gnd cell_6t
Xbit_r105_c39 bl_39 br_39 wl_105 vdd gnd cell_6t
Xbit_r106_c39 bl_39 br_39 wl_106 vdd gnd cell_6t
Xbit_r107_c39 bl_39 br_39 wl_107 vdd gnd cell_6t
Xbit_r108_c39 bl_39 br_39 wl_108 vdd gnd cell_6t
Xbit_r109_c39 bl_39 br_39 wl_109 vdd gnd cell_6t
Xbit_r110_c39 bl_39 br_39 wl_110 vdd gnd cell_6t
Xbit_r111_c39 bl_39 br_39 wl_111 vdd gnd cell_6t
Xbit_r112_c39 bl_39 br_39 wl_112 vdd gnd cell_6t
Xbit_r113_c39 bl_39 br_39 wl_113 vdd gnd cell_6t
Xbit_r114_c39 bl_39 br_39 wl_114 vdd gnd cell_6t
Xbit_r115_c39 bl_39 br_39 wl_115 vdd gnd cell_6t
Xbit_r116_c39 bl_39 br_39 wl_116 vdd gnd cell_6t
Xbit_r117_c39 bl_39 br_39 wl_117 vdd gnd cell_6t
Xbit_r118_c39 bl_39 br_39 wl_118 vdd gnd cell_6t
Xbit_r119_c39 bl_39 br_39 wl_119 vdd gnd cell_6t
Xbit_r120_c39 bl_39 br_39 wl_120 vdd gnd cell_6t
Xbit_r121_c39 bl_39 br_39 wl_121 vdd gnd cell_6t
Xbit_r122_c39 bl_39 br_39 wl_122 vdd gnd cell_6t
Xbit_r123_c39 bl_39 br_39 wl_123 vdd gnd cell_6t
Xbit_r124_c39 bl_39 br_39 wl_124 vdd gnd cell_6t
Xbit_r125_c39 bl_39 br_39 wl_125 vdd gnd cell_6t
Xbit_r126_c39 bl_39 br_39 wl_126 vdd gnd cell_6t
Xbit_r127_c39 bl_39 br_39 wl_127 vdd gnd cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd cell_6t
Xbit_r1_c40 bl_40 br_40 wl_1 vdd gnd cell_6t
Xbit_r2_c40 bl_40 br_40 wl_2 vdd gnd cell_6t
Xbit_r3_c40 bl_40 br_40 wl_3 vdd gnd cell_6t
Xbit_r4_c40 bl_40 br_40 wl_4 vdd gnd cell_6t
Xbit_r5_c40 bl_40 br_40 wl_5 vdd gnd cell_6t
Xbit_r6_c40 bl_40 br_40 wl_6 vdd gnd cell_6t
Xbit_r7_c40 bl_40 br_40 wl_7 vdd gnd cell_6t
Xbit_r8_c40 bl_40 br_40 wl_8 vdd gnd cell_6t
Xbit_r9_c40 bl_40 br_40 wl_9 vdd gnd cell_6t
Xbit_r10_c40 bl_40 br_40 wl_10 vdd gnd cell_6t
Xbit_r11_c40 bl_40 br_40 wl_11 vdd gnd cell_6t
Xbit_r12_c40 bl_40 br_40 wl_12 vdd gnd cell_6t
Xbit_r13_c40 bl_40 br_40 wl_13 vdd gnd cell_6t
Xbit_r14_c40 bl_40 br_40 wl_14 vdd gnd cell_6t
Xbit_r15_c40 bl_40 br_40 wl_15 vdd gnd cell_6t
Xbit_r16_c40 bl_40 br_40 wl_16 vdd gnd cell_6t
Xbit_r17_c40 bl_40 br_40 wl_17 vdd gnd cell_6t
Xbit_r18_c40 bl_40 br_40 wl_18 vdd gnd cell_6t
Xbit_r19_c40 bl_40 br_40 wl_19 vdd gnd cell_6t
Xbit_r20_c40 bl_40 br_40 wl_20 vdd gnd cell_6t
Xbit_r21_c40 bl_40 br_40 wl_21 vdd gnd cell_6t
Xbit_r22_c40 bl_40 br_40 wl_22 vdd gnd cell_6t
Xbit_r23_c40 bl_40 br_40 wl_23 vdd gnd cell_6t
Xbit_r24_c40 bl_40 br_40 wl_24 vdd gnd cell_6t
Xbit_r25_c40 bl_40 br_40 wl_25 vdd gnd cell_6t
Xbit_r26_c40 bl_40 br_40 wl_26 vdd gnd cell_6t
Xbit_r27_c40 bl_40 br_40 wl_27 vdd gnd cell_6t
Xbit_r28_c40 bl_40 br_40 wl_28 vdd gnd cell_6t
Xbit_r29_c40 bl_40 br_40 wl_29 vdd gnd cell_6t
Xbit_r30_c40 bl_40 br_40 wl_30 vdd gnd cell_6t
Xbit_r31_c40 bl_40 br_40 wl_31 vdd gnd cell_6t
Xbit_r32_c40 bl_40 br_40 wl_32 vdd gnd cell_6t
Xbit_r33_c40 bl_40 br_40 wl_33 vdd gnd cell_6t
Xbit_r34_c40 bl_40 br_40 wl_34 vdd gnd cell_6t
Xbit_r35_c40 bl_40 br_40 wl_35 vdd gnd cell_6t
Xbit_r36_c40 bl_40 br_40 wl_36 vdd gnd cell_6t
Xbit_r37_c40 bl_40 br_40 wl_37 vdd gnd cell_6t
Xbit_r38_c40 bl_40 br_40 wl_38 vdd gnd cell_6t
Xbit_r39_c40 bl_40 br_40 wl_39 vdd gnd cell_6t
Xbit_r40_c40 bl_40 br_40 wl_40 vdd gnd cell_6t
Xbit_r41_c40 bl_40 br_40 wl_41 vdd gnd cell_6t
Xbit_r42_c40 bl_40 br_40 wl_42 vdd gnd cell_6t
Xbit_r43_c40 bl_40 br_40 wl_43 vdd gnd cell_6t
Xbit_r44_c40 bl_40 br_40 wl_44 vdd gnd cell_6t
Xbit_r45_c40 bl_40 br_40 wl_45 vdd gnd cell_6t
Xbit_r46_c40 bl_40 br_40 wl_46 vdd gnd cell_6t
Xbit_r47_c40 bl_40 br_40 wl_47 vdd gnd cell_6t
Xbit_r48_c40 bl_40 br_40 wl_48 vdd gnd cell_6t
Xbit_r49_c40 bl_40 br_40 wl_49 vdd gnd cell_6t
Xbit_r50_c40 bl_40 br_40 wl_50 vdd gnd cell_6t
Xbit_r51_c40 bl_40 br_40 wl_51 vdd gnd cell_6t
Xbit_r52_c40 bl_40 br_40 wl_52 vdd gnd cell_6t
Xbit_r53_c40 bl_40 br_40 wl_53 vdd gnd cell_6t
Xbit_r54_c40 bl_40 br_40 wl_54 vdd gnd cell_6t
Xbit_r55_c40 bl_40 br_40 wl_55 vdd gnd cell_6t
Xbit_r56_c40 bl_40 br_40 wl_56 vdd gnd cell_6t
Xbit_r57_c40 bl_40 br_40 wl_57 vdd gnd cell_6t
Xbit_r58_c40 bl_40 br_40 wl_58 vdd gnd cell_6t
Xbit_r59_c40 bl_40 br_40 wl_59 vdd gnd cell_6t
Xbit_r60_c40 bl_40 br_40 wl_60 vdd gnd cell_6t
Xbit_r61_c40 bl_40 br_40 wl_61 vdd gnd cell_6t
Xbit_r62_c40 bl_40 br_40 wl_62 vdd gnd cell_6t
Xbit_r63_c40 bl_40 br_40 wl_63 vdd gnd cell_6t
Xbit_r64_c40 bl_40 br_40 wl_64 vdd gnd cell_6t
Xbit_r65_c40 bl_40 br_40 wl_65 vdd gnd cell_6t
Xbit_r66_c40 bl_40 br_40 wl_66 vdd gnd cell_6t
Xbit_r67_c40 bl_40 br_40 wl_67 vdd gnd cell_6t
Xbit_r68_c40 bl_40 br_40 wl_68 vdd gnd cell_6t
Xbit_r69_c40 bl_40 br_40 wl_69 vdd gnd cell_6t
Xbit_r70_c40 bl_40 br_40 wl_70 vdd gnd cell_6t
Xbit_r71_c40 bl_40 br_40 wl_71 vdd gnd cell_6t
Xbit_r72_c40 bl_40 br_40 wl_72 vdd gnd cell_6t
Xbit_r73_c40 bl_40 br_40 wl_73 vdd gnd cell_6t
Xbit_r74_c40 bl_40 br_40 wl_74 vdd gnd cell_6t
Xbit_r75_c40 bl_40 br_40 wl_75 vdd gnd cell_6t
Xbit_r76_c40 bl_40 br_40 wl_76 vdd gnd cell_6t
Xbit_r77_c40 bl_40 br_40 wl_77 vdd gnd cell_6t
Xbit_r78_c40 bl_40 br_40 wl_78 vdd gnd cell_6t
Xbit_r79_c40 bl_40 br_40 wl_79 vdd gnd cell_6t
Xbit_r80_c40 bl_40 br_40 wl_80 vdd gnd cell_6t
Xbit_r81_c40 bl_40 br_40 wl_81 vdd gnd cell_6t
Xbit_r82_c40 bl_40 br_40 wl_82 vdd gnd cell_6t
Xbit_r83_c40 bl_40 br_40 wl_83 vdd gnd cell_6t
Xbit_r84_c40 bl_40 br_40 wl_84 vdd gnd cell_6t
Xbit_r85_c40 bl_40 br_40 wl_85 vdd gnd cell_6t
Xbit_r86_c40 bl_40 br_40 wl_86 vdd gnd cell_6t
Xbit_r87_c40 bl_40 br_40 wl_87 vdd gnd cell_6t
Xbit_r88_c40 bl_40 br_40 wl_88 vdd gnd cell_6t
Xbit_r89_c40 bl_40 br_40 wl_89 vdd gnd cell_6t
Xbit_r90_c40 bl_40 br_40 wl_90 vdd gnd cell_6t
Xbit_r91_c40 bl_40 br_40 wl_91 vdd gnd cell_6t
Xbit_r92_c40 bl_40 br_40 wl_92 vdd gnd cell_6t
Xbit_r93_c40 bl_40 br_40 wl_93 vdd gnd cell_6t
Xbit_r94_c40 bl_40 br_40 wl_94 vdd gnd cell_6t
Xbit_r95_c40 bl_40 br_40 wl_95 vdd gnd cell_6t
Xbit_r96_c40 bl_40 br_40 wl_96 vdd gnd cell_6t
Xbit_r97_c40 bl_40 br_40 wl_97 vdd gnd cell_6t
Xbit_r98_c40 bl_40 br_40 wl_98 vdd gnd cell_6t
Xbit_r99_c40 bl_40 br_40 wl_99 vdd gnd cell_6t
Xbit_r100_c40 bl_40 br_40 wl_100 vdd gnd cell_6t
Xbit_r101_c40 bl_40 br_40 wl_101 vdd gnd cell_6t
Xbit_r102_c40 bl_40 br_40 wl_102 vdd gnd cell_6t
Xbit_r103_c40 bl_40 br_40 wl_103 vdd gnd cell_6t
Xbit_r104_c40 bl_40 br_40 wl_104 vdd gnd cell_6t
Xbit_r105_c40 bl_40 br_40 wl_105 vdd gnd cell_6t
Xbit_r106_c40 bl_40 br_40 wl_106 vdd gnd cell_6t
Xbit_r107_c40 bl_40 br_40 wl_107 vdd gnd cell_6t
Xbit_r108_c40 bl_40 br_40 wl_108 vdd gnd cell_6t
Xbit_r109_c40 bl_40 br_40 wl_109 vdd gnd cell_6t
Xbit_r110_c40 bl_40 br_40 wl_110 vdd gnd cell_6t
Xbit_r111_c40 bl_40 br_40 wl_111 vdd gnd cell_6t
Xbit_r112_c40 bl_40 br_40 wl_112 vdd gnd cell_6t
Xbit_r113_c40 bl_40 br_40 wl_113 vdd gnd cell_6t
Xbit_r114_c40 bl_40 br_40 wl_114 vdd gnd cell_6t
Xbit_r115_c40 bl_40 br_40 wl_115 vdd gnd cell_6t
Xbit_r116_c40 bl_40 br_40 wl_116 vdd gnd cell_6t
Xbit_r117_c40 bl_40 br_40 wl_117 vdd gnd cell_6t
Xbit_r118_c40 bl_40 br_40 wl_118 vdd gnd cell_6t
Xbit_r119_c40 bl_40 br_40 wl_119 vdd gnd cell_6t
Xbit_r120_c40 bl_40 br_40 wl_120 vdd gnd cell_6t
Xbit_r121_c40 bl_40 br_40 wl_121 vdd gnd cell_6t
Xbit_r122_c40 bl_40 br_40 wl_122 vdd gnd cell_6t
Xbit_r123_c40 bl_40 br_40 wl_123 vdd gnd cell_6t
Xbit_r124_c40 bl_40 br_40 wl_124 vdd gnd cell_6t
Xbit_r125_c40 bl_40 br_40 wl_125 vdd gnd cell_6t
Xbit_r126_c40 bl_40 br_40 wl_126 vdd gnd cell_6t
Xbit_r127_c40 bl_40 br_40 wl_127 vdd gnd cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd cell_6t
Xbit_r1_c41 bl_41 br_41 wl_1 vdd gnd cell_6t
Xbit_r2_c41 bl_41 br_41 wl_2 vdd gnd cell_6t
Xbit_r3_c41 bl_41 br_41 wl_3 vdd gnd cell_6t
Xbit_r4_c41 bl_41 br_41 wl_4 vdd gnd cell_6t
Xbit_r5_c41 bl_41 br_41 wl_5 vdd gnd cell_6t
Xbit_r6_c41 bl_41 br_41 wl_6 vdd gnd cell_6t
Xbit_r7_c41 bl_41 br_41 wl_7 vdd gnd cell_6t
Xbit_r8_c41 bl_41 br_41 wl_8 vdd gnd cell_6t
Xbit_r9_c41 bl_41 br_41 wl_9 vdd gnd cell_6t
Xbit_r10_c41 bl_41 br_41 wl_10 vdd gnd cell_6t
Xbit_r11_c41 bl_41 br_41 wl_11 vdd gnd cell_6t
Xbit_r12_c41 bl_41 br_41 wl_12 vdd gnd cell_6t
Xbit_r13_c41 bl_41 br_41 wl_13 vdd gnd cell_6t
Xbit_r14_c41 bl_41 br_41 wl_14 vdd gnd cell_6t
Xbit_r15_c41 bl_41 br_41 wl_15 vdd gnd cell_6t
Xbit_r16_c41 bl_41 br_41 wl_16 vdd gnd cell_6t
Xbit_r17_c41 bl_41 br_41 wl_17 vdd gnd cell_6t
Xbit_r18_c41 bl_41 br_41 wl_18 vdd gnd cell_6t
Xbit_r19_c41 bl_41 br_41 wl_19 vdd gnd cell_6t
Xbit_r20_c41 bl_41 br_41 wl_20 vdd gnd cell_6t
Xbit_r21_c41 bl_41 br_41 wl_21 vdd gnd cell_6t
Xbit_r22_c41 bl_41 br_41 wl_22 vdd gnd cell_6t
Xbit_r23_c41 bl_41 br_41 wl_23 vdd gnd cell_6t
Xbit_r24_c41 bl_41 br_41 wl_24 vdd gnd cell_6t
Xbit_r25_c41 bl_41 br_41 wl_25 vdd gnd cell_6t
Xbit_r26_c41 bl_41 br_41 wl_26 vdd gnd cell_6t
Xbit_r27_c41 bl_41 br_41 wl_27 vdd gnd cell_6t
Xbit_r28_c41 bl_41 br_41 wl_28 vdd gnd cell_6t
Xbit_r29_c41 bl_41 br_41 wl_29 vdd gnd cell_6t
Xbit_r30_c41 bl_41 br_41 wl_30 vdd gnd cell_6t
Xbit_r31_c41 bl_41 br_41 wl_31 vdd gnd cell_6t
Xbit_r32_c41 bl_41 br_41 wl_32 vdd gnd cell_6t
Xbit_r33_c41 bl_41 br_41 wl_33 vdd gnd cell_6t
Xbit_r34_c41 bl_41 br_41 wl_34 vdd gnd cell_6t
Xbit_r35_c41 bl_41 br_41 wl_35 vdd gnd cell_6t
Xbit_r36_c41 bl_41 br_41 wl_36 vdd gnd cell_6t
Xbit_r37_c41 bl_41 br_41 wl_37 vdd gnd cell_6t
Xbit_r38_c41 bl_41 br_41 wl_38 vdd gnd cell_6t
Xbit_r39_c41 bl_41 br_41 wl_39 vdd gnd cell_6t
Xbit_r40_c41 bl_41 br_41 wl_40 vdd gnd cell_6t
Xbit_r41_c41 bl_41 br_41 wl_41 vdd gnd cell_6t
Xbit_r42_c41 bl_41 br_41 wl_42 vdd gnd cell_6t
Xbit_r43_c41 bl_41 br_41 wl_43 vdd gnd cell_6t
Xbit_r44_c41 bl_41 br_41 wl_44 vdd gnd cell_6t
Xbit_r45_c41 bl_41 br_41 wl_45 vdd gnd cell_6t
Xbit_r46_c41 bl_41 br_41 wl_46 vdd gnd cell_6t
Xbit_r47_c41 bl_41 br_41 wl_47 vdd gnd cell_6t
Xbit_r48_c41 bl_41 br_41 wl_48 vdd gnd cell_6t
Xbit_r49_c41 bl_41 br_41 wl_49 vdd gnd cell_6t
Xbit_r50_c41 bl_41 br_41 wl_50 vdd gnd cell_6t
Xbit_r51_c41 bl_41 br_41 wl_51 vdd gnd cell_6t
Xbit_r52_c41 bl_41 br_41 wl_52 vdd gnd cell_6t
Xbit_r53_c41 bl_41 br_41 wl_53 vdd gnd cell_6t
Xbit_r54_c41 bl_41 br_41 wl_54 vdd gnd cell_6t
Xbit_r55_c41 bl_41 br_41 wl_55 vdd gnd cell_6t
Xbit_r56_c41 bl_41 br_41 wl_56 vdd gnd cell_6t
Xbit_r57_c41 bl_41 br_41 wl_57 vdd gnd cell_6t
Xbit_r58_c41 bl_41 br_41 wl_58 vdd gnd cell_6t
Xbit_r59_c41 bl_41 br_41 wl_59 vdd gnd cell_6t
Xbit_r60_c41 bl_41 br_41 wl_60 vdd gnd cell_6t
Xbit_r61_c41 bl_41 br_41 wl_61 vdd gnd cell_6t
Xbit_r62_c41 bl_41 br_41 wl_62 vdd gnd cell_6t
Xbit_r63_c41 bl_41 br_41 wl_63 vdd gnd cell_6t
Xbit_r64_c41 bl_41 br_41 wl_64 vdd gnd cell_6t
Xbit_r65_c41 bl_41 br_41 wl_65 vdd gnd cell_6t
Xbit_r66_c41 bl_41 br_41 wl_66 vdd gnd cell_6t
Xbit_r67_c41 bl_41 br_41 wl_67 vdd gnd cell_6t
Xbit_r68_c41 bl_41 br_41 wl_68 vdd gnd cell_6t
Xbit_r69_c41 bl_41 br_41 wl_69 vdd gnd cell_6t
Xbit_r70_c41 bl_41 br_41 wl_70 vdd gnd cell_6t
Xbit_r71_c41 bl_41 br_41 wl_71 vdd gnd cell_6t
Xbit_r72_c41 bl_41 br_41 wl_72 vdd gnd cell_6t
Xbit_r73_c41 bl_41 br_41 wl_73 vdd gnd cell_6t
Xbit_r74_c41 bl_41 br_41 wl_74 vdd gnd cell_6t
Xbit_r75_c41 bl_41 br_41 wl_75 vdd gnd cell_6t
Xbit_r76_c41 bl_41 br_41 wl_76 vdd gnd cell_6t
Xbit_r77_c41 bl_41 br_41 wl_77 vdd gnd cell_6t
Xbit_r78_c41 bl_41 br_41 wl_78 vdd gnd cell_6t
Xbit_r79_c41 bl_41 br_41 wl_79 vdd gnd cell_6t
Xbit_r80_c41 bl_41 br_41 wl_80 vdd gnd cell_6t
Xbit_r81_c41 bl_41 br_41 wl_81 vdd gnd cell_6t
Xbit_r82_c41 bl_41 br_41 wl_82 vdd gnd cell_6t
Xbit_r83_c41 bl_41 br_41 wl_83 vdd gnd cell_6t
Xbit_r84_c41 bl_41 br_41 wl_84 vdd gnd cell_6t
Xbit_r85_c41 bl_41 br_41 wl_85 vdd gnd cell_6t
Xbit_r86_c41 bl_41 br_41 wl_86 vdd gnd cell_6t
Xbit_r87_c41 bl_41 br_41 wl_87 vdd gnd cell_6t
Xbit_r88_c41 bl_41 br_41 wl_88 vdd gnd cell_6t
Xbit_r89_c41 bl_41 br_41 wl_89 vdd gnd cell_6t
Xbit_r90_c41 bl_41 br_41 wl_90 vdd gnd cell_6t
Xbit_r91_c41 bl_41 br_41 wl_91 vdd gnd cell_6t
Xbit_r92_c41 bl_41 br_41 wl_92 vdd gnd cell_6t
Xbit_r93_c41 bl_41 br_41 wl_93 vdd gnd cell_6t
Xbit_r94_c41 bl_41 br_41 wl_94 vdd gnd cell_6t
Xbit_r95_c41 bl_41 br_41 wl_95 vdd gnd cell_6t
Xbit_r96_c41 bl_41 br_41 wl_96 vdd gnd cell_6t
Xbit_r97_c41 bl_41 br_41 wl_97 vdd gnd cell_6t
Xbit_r98_c41 bl_41 br_41 wl_98 vdd gnd cell_6t
Xbit_r99_c41 bl_41 br_41 wl_99 vdd gnd cell_6t
Xbit_r100_c41 bl_41 br_41 wl_100 vdd gnd cell_6t
Xbit_r101_c41 bl_41 br_41 wl_101 vdd gnd cell_6t
Xbit_r102_c41 bl_41 br_41 wl_102 vdd gnd cell_6t
Xbit_r103_c41 bl_41 br_41 wl_103 vdd gnd cell_6t
Xbit_r104_c41 bl_41 br_41 wl_104 vdd gnd cell_6t
Xbit_r105_c41 bl_41 br_41 wl_105 vdd gnd cell_6t
Xbit_r106_c41 bl_41 br_41 wl_106 vdd gnd cell_6t
Xbit_r107_c41 bl_41 br_41 wl_107 vdd gnd cell_6t
Xbit_r108_c41 bl_41 br_41 wl_108 vdd gnd cell_6t
Xbit_r109_c41 bl_41 br_41 wl_109 vdd gnd cell_6t
Xbit_r110_c41 bl_41 br_41 wl_110 vdd gnd cell_6t
Xbit_r111_c41 bl_41 br_41 wl_111 vdd gnd cell_6t
Xbit_r112_c41 bl_41 br_41 wl_112 vdd gnd cell_6t
Xbit_r113_c41 bl_41 br_41 wl_113 vdd gnd cell_6t
Xbit_r114_c41 bl_41 br_41 wl_114 vdd gnd cell_6t
Xbit_r115_c41 bl_41 br_41 wl_115 vdd gnd cell_6t
Xbit_r116_c41 bl_41 br_41 wl_116 vdd gnd cell_6t
Xbit_r117_c41 bl_41 br_41 wl_117 vdd gnd cell_6t
Xbit_r118_c41 bl_41 br_41 wl_118 vdd gnd cell_6t
Xbit_r119_c41 bl_41 br_41 wl_119 vdd gnd cell_6t
Xbit_r120_c41 bl_41 br_41 wl_120 vdd gnd cell_6t
Xbit_r121_c41 bl_41 br_41 wl_121 vdd gnd cell_6t
Xbit_r122_c41 bl_41 br_41 wl_122 vdd gnd cell_6t
Xbit_r123_c41 bl_41 br_41 wl_123 vdd gnd cell_6t
Xbit_r124_c41 bl_41 br_41 wl_124 vdd gnd cell_6t
Xbit_r125_c41 bl_41 br_41 wl_125 vdd gnd cell_6t
Xbit_r126_c41 bl_41 br_41 wl_126 vdd gnd cell_6t
Xbit_r127_c41 bl_41 br_41 wl_127 vdd gnd cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd cell_6t
Xbit_r1_c42 bl_42 br_42 wl_1 vdd gnd cell_6t
Xbit_r2_c42 bl_42 br_42 wl_2 vdd gnd cell_6t
Xbit_r3_c42 bl_42 br_42 wl_3 vdd gnd cell_6t
Xbit_r4_c42 bl_42 br_42 wl_4 vdd gnd cell_6t
Xbit_r5_c42 bl_42 br_42 wl_5 vdd gnd cell_6t
Xbit_r6_c42 bl_42 br_42 wl_6 vdd gnd cell_6t
Xbit_r7_c42 bl_42 br_42 wl_7 vdd gnd cell_6t
Xbit_r8_c42 bl_42 br_42 wl_8 vdd gnd cell_6t
Xbit_r9_c42 bl_42 br_42 wl_9 vdd gnd cell_6t
Xbit_r10_c42 bl_42 br_42 wl_10 vdd gnd cell_6t
Xbit_r11_c42 bl_42 br_42 wl_11 vdd gnd cell_6t
Xbit_r12_c42 bl_42 br_42 wl_12 vdd gnd cell_6t
Xbit_r13_c42 bl_42 br_42 wl_13 vdd gnd cell_6t
Xbit_r14_c42 bl_42 br_42 wl_14 vdd gnd cell_6t
Xbit_r15_c42 bl_42 br_42 wl_15 vdd gnd cell_6t
Xbit_r16_c42 bl_42 br_42 wl_16 vdd gnd cell_6t
Xbit_r17_c42 bl_42 br_42 wl_17 vdd gnd cell_6t
Xbit_r18_c42 bl_42 br_42 wl_18 vdd gnd cell_6t
Xbit_r19_c42 bl_42 br_42 wl_19 vdd gnd cell_6t
Xbit_r20_c42 bl_42 br_42 wl_20 vdd gnd cell_6t
Xbit_r21_c42 bl_42 br_42 wl_21 vdd gnd cell_6t
Xbit_r22_c42 bl_42 br_42 wl_22 vdd gnd cell_6t
Xbit_r23_c42 bl_42 br_42 wl_23 vdd gnd cell_6t
Xbit_r24_c42 bl_42 br_42 wl_24 vdd gnd cell_6t
Xbit_r25_c42 bl_42 br_42 wl_25 vdd gnd cell_6t
Xbit_r26_c42 bl_42 br_42 wl_26 vdd gnd cell_6t
Xbit_r27_c42 bl_42 br_42 wl_27 vdd gnd cell_6t
Xbit_r28_c42 bl_42 br_42 wl_28 vdd gnd cell_6t
Xbit_r29_c42 bl_42 br_42 wl_29 vdd gnd cell_6t
Xbit_r30_c42 bl_42 br_42 wl_30 vdd gnd cell_6t
Xbit_r31_c42 bl_42 br_42 wl_31 vdd gnd cell_6t
Xbit_r32_c42 bl_42 br_42 wl_32 vdd gnd cell_6t
Xbit_r33_c42 bl_42 br_42 wl_33 vdd gnd cell_6t
Xbit_r34_c42 bl_42 br_42 wl_34 vdd gnd cell_6t
Xbit_r35_c42 bl_42 br_42 wl_35 vdd gnd cell_6t
Xbit_r36_c42 bl_42 br_42 wl_36 vdd gnd cell_6t
Xbit_r37_c42 bl_42 br_42 wl_37 vdd gnd cell_6t
Xbit_r38_c42 bl_42 br_42 wl_38 vdd gnd cell_6t
Xbit_r39_c42 bl_42 br_42 wl_39 vdd gnd cell_6t
Xbit_r40_c42 bl_42 br_42 wl_40 vdd gnd cell_6t
Xbit_r41_c42 bl_42 br_42 wl_41 vdd gnd cell_6t
Xbit_r42_c42 bl_42 br_42 wl_42 vdd gnd cell_6t
Xbit_r43_c42 bl_42 br_42 wl_43 vdd gnd cell_6t
Xbit_r44_c42 bl_42 br_42 wl_44 vdd gnd cell_6t
Xbit_r45_c42 bl_42 br_42 wl_45 vdd gnd cell_6t
Xbit_r46_c42 bl_42 br_42 wl_46 vdd gnd cell_6t
Xbit_r47_c42 bl_42 br_42 wl_47 vdd gnd cell_6t
Xbit_r48_c42 bl_42 br_42 wl_48 vdd gnd cell_6t
Xbit_r49_c42 bl_42 br_42 wl_49 vdd gnd cell_6t
Xbit_r50_c42 bl_42 br_42 wl_50 vdd gnd cell_6t
Xbit_r51_c42 bl_42 br_42 wl_51 vdd gnd cell_6t
Xbit_r52_c42 bl_42 br_42 wl_52 vdd gnd cell_6t
Xbit_r53_c42 bl_42 br_42 wl_53 vdd gnd cell_6t
Xbit_r54_c42 bl_42 br_42 wl_54 vdd gnd cell_6t
Xbit_r55_c42 bl_42 br_42 wl_55 vdd gnd cell_6t
Xbit_r56_c42 bl_42 br_42 wl_56 vdd gnd cell_6t
Xbit_r57_c42 bl_42 br_42 wl_57 vdd gnd cell_6t
Xbit_r58_c42 bl_42 br_42 wl_58 vdd gnd cell_6t
Xbit_r59_c42 bl_42 br_42 wl_59 vdd gnd cell_6t
Xbit_r60_c42 bl_42 br_42 wl_60 vdd gnd cell_6t
Xbit_r61_c42 bl_42 br_42 wl_61 vdd gnd cell_6t
Xbit_r62_c42 bl_42 br_42 wl_62 vdd gnd cell_6t
Xbit_r63_c42 bl_42 br_42 wl_63 vdd gnd cell_6t
Xbit_r64_c42 bl_42 br_42 wl_64 vdd gnd cell_6t
Xbit_r65_c42 bl_42 br_42 wl_65 vdd gnd cell_6t
Xbit_r66_c42 bl_42 br_42 wl_66 vdd gnd cell_6t
Xbit_r67_c42 bl_42 br_42 wl_67 vdd gnd cell_6t
Xbit_r68_c42 bl_42 br_42 wl_68 vdd gnd cell_6t
Xbit_r69_c42 bl_42 br_42 wl_69 vdd gnd cell_6t
Xbit_r70_c42 bl_42 br_42 wl_70 vdd gnd cell_6t
Xbit_r71_c42 bl_42 br_42 wl_71 vdd gnd cell_6t
Xbit_r72_c42 bl_42 br_42 wl_72 vdd gnd cell_6t
Xbit_r73_c42 bl_42 br_42 wl_73 vdd gnd cell_6t
Xbit_r74_c42 bl_42 br_42 wl_74 vdd gnd cell_6t
Xbit_r75_c42 bl_42 br_42 wl_75 vdd gnd cell_6t
Xbit_r76_c42 bl_42 br_42 wl_76 vdd gnd cell_6t
Xbit_r77_c42 bl_42 br_42 wl_77 vdd gnd cell_6t
Xbit_r78_c42 bl_42 br_42 wl_78 vdd gnd cell_6t
Xbit_r79_c42 bl_42 br_42 wl_79 vdd gnd cell_6t
Xbit_r80_c42 bl_42 br_42 wl_80 vdd gnd cell_6t
Xbit_r81_c42 bl_42 br_42 wl_81 vdd gnd cell_6t
Xbit_r82_c42 bl_42 br_42 wl_82 vdd gnd cell_6t
Xbit_r83_c42 bl_42 br_42 wl_83 vdd gnd cell_6t
Xbit_r84_c42 bl_42 br_42 wl_84 vdd gnd cell_6t
Xbit_r85_c42 bl_42 br_42 wl_85 vdd gnd cell_6t
Xbit_r86_c42 bl_42 br_42 wl_86 vdd gnd cell_6t
Xbit_r87_c42 bl_42 br_42 wl_87 vdd gnd cell_6t
Xbit_r88_c42 bl_42 br_42 wl_88 vdd gnd cell_6t
Xbit_r89_c42 bl_42 br_42 wl_89 vdd gnd cell_6t
Xbit_r90_c42 bl_42 br_42 wl_90 vdd gnd cell_6t
Xbit_r91_c42 bl_42 br_42 wl_91 vdd gnd cell_6t
Xbit_r92_c42 bl_42 br_42 wl_92 vdd gnd cell_6t
Xbit_r93_c42 bl_42 br_42 wl_93 vdd gnd cell_6t
Xbit_r94_c42 bl_42 br_42 wl_94 vdd gnd cell_6t
Xbit_r95_c42 bl_42 br_42 wl_95 vdd gnd cell_6t
Xbit_r96_c42 bl_42 br_42 wl_96 vdd gnd cell_6t
Xbit_r97_c42 bl_42 br_42 wl_97 vdd gnd cell_6t
Xbit_r98_c42 bl_42 br_42 wl_98 vdd gnd cell_6t
Xbit_r99_c42 bl_42 br_42 wl_99 vdd gnd cell_6t
Xbit_r100_c42 bl_42 br_42 wl_100 vdd gnd cell_6t
Xbit_r101_c42 bl_42 br_42 wl_101 vdd gnd cell_6t
Xbit_r102_c42 bl_42 br_42 wl_102 vdd gnd cell_6t
Xbit_r103_c42 bl_42 br_42 wl_103 vdd gnd cell_6t
Xbit_r104_c42 bl_42 br_42 wl_104 vdd gnd cell_6t
Xbit_r105_c42 bl_42 br_42 wl_105 vdd gnd cell_6t
Xbit_r106_c42 bl_42 br_42 wl_106 vdd gnd cell_6t
Xbit_r107_c42 bl_42 br_42 wl_107 vdd gnd cell_6t
Xbit_r108_c42 bl_42 br_42 wl_108 vdd gnd cell_6t
Xbit_r109_c42 bl_42 br_42 wl_109 vdd gnd cell_6t
Xbit_r110_c42 bl_42 br_42 wl_110 vdd gnd cell_6t
Xbit_r111_c42 bl_42 br_42 wl_111 vdd gnd cell_6t
Xbit_r112_c42 bl_42 br_42 wl_112 vdd gnd cell_6t
Xbit_r113_c42 bl_42 br_42 wl_113 vdd gnd cell_6t
Xbit_r114_c42 bl_42 br_42 wl_114 vdd gnd cell_6t
Xbit_r115_c42 bl_42 br_42 wl_115 vdd gnd cell_6t
Xbit_r116_c42 bl_42 br_42 wl_116 vdd gnd cell_6t
Xbit_r117_c42 bl_42 br_42 wl_117 vdd gnd cell_6t
Xbit_r118_c42 bl_42 br_42 wl_118 vdd gnd cell_6t
Xbit_r119_c42 bl_42 br_42 wl_119 vdd gnd cell_6t
Xbit_r120_c42 bl_42 br_42 wl_120 vdd gnd cell_6t
Xbit_r121_c42 bl_42 br_42 wl_121 vdd gnd cell_6t
Xbit_r122_c42 bl_42 br_42 wl_122 vdd gnd cell_6t
Xbit_r123_c42 bl_42 br_42 wl_123 vdd gnd cell_6t
Xbit_r124_c42 bl_42 br_42 wl_124 vdd gnd cell_6t
Xbit_r125_c42 bl_42 br_42 wl_125 vdd gnd cell_6t
Xbit_r126_c42 bl_42 br_42 wl_126 vdd gnd cell_6t
Xbit_r127_c42 bl_42 br_42 wl_127 vdd gnd cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd cell_6t
Xbit_r1_c43 bl_43 br_43 wl_1 vdd gnd cell_6t
Xbit_r2_c43 bl_43 br_43 wl_2 vdd gnd cell_6t
Xbit_r3_c43 bl_43 br_43 wl_3 vdd gnd cell_6t
Xbit_r4_c43 bl_43 br_43 wl_4 vdd gnd cell_6t
Xbit_r5_c43 bl_43 br_43 wl_5 vdd gnd cell_6t
Xbit_r6_c43 bl_43 br_43 wl_6 vdd gnd cell_6t
Xbit_r7_c43 bl_43 br_43 wl_7 vdd gnd cell_6t
Xbit_r8_c43 bl_43 br_43 wl_8 vdd gnd cell_6t
Xbit_r9_c43 bl_43 br_43 wl_9 vdd gnd cell_6t
Xbit_r10_c43 bl_43 br_43 wl_10 vdd gnd cell_6t
Xbit_r11_c43 bl_43 br_43 wl_11 vdd gnd cell_6t
Xbit_r12_c43 bl_43 br_43 wl_12 vdd gnd cell_6t
Xbit_r13_c43 bl_43 br_43 wl_13 vdd gnd cell_6t
Xbit_r14_c43 bl_43 br_43 wl_14 vdd gnd cell_6t
Xbit_r15_c43 bl_43 br_43 wl_15 vdd gnd cell_6t
Xbit_r16_c43 bl_43 br_43 wl_16 vdd gnd cell_6t
Xbit_r17_c43 bl_43 br_43 wl_17 vdd gnd cell_6t
Xbit_r18_c43 bl_43 br_43 wl_18 vdd gnd cell_6t
Xbit_r19_c43 bl_43 br_43 wl_19 vdd gnd cell_6t
Xbit_r20_c43 bl_43 br_43 wl_20 vdd gnd cell_6t
Xbit_r21_c43 bl_43 br_43 wl_21 vdd gnd cell_6t
Xbit_r22_c43 bl_43 br_43 wl_22 vdd gnd cell_6t
Xbit_r23_c43 bl_43 br_43 wl_23 vdd gnd cell_6t
Xbit_r24_c43 bl_43 br_43 wl_24 vdd gnd cell_6t
Xbit_r25_c43 bl_43 br_43 wl_25 vdd gnd cell_6t
Xbit_r26_c43 bl_43 br_43 wl_26 vdd gnd cell_6t
Xbit_r27_c43 bl_43 br_43 wl_27 vdd gnd cell_6t
Xbit_r28_c43 bl_43 br_43 wl_28 vdd gnd cell_6t
Xbit_r29_c43 bl_43 br_43 wl_29 vdd gnd cell_6t
Xbit_r30_c43 bl_43 br_43 wl_30 vdd gnd cell_6t
Xbit_r31_c43 bl_43 br_43 wl_31 vdd gnd cell_6t
Xbit_r32_c43 bl_43 br_43 wl_32 vdd gnd cell_6t
Xbit_r33_c43 bl_43 br_43 wl_33 vdd gnd cell_6t
Xbit_r34_c43 bl_43 br_43 wl_34 vdd gnd cell_6t
Xbit_r35_c43 bl_43 br_43 wl_35 vdd gnd cell_6t
Xbit_r36_c43 bl_43 br_43 wl_36 vdd gnd cell_6t
Xbit_r37_c43 bl_43 br_43 wl_37 vdd gnd cell_6t
Xbit_r38_c43 bl_43 br_43 wl_38 vdd gnd cell_6t
Xbit_r39_c43 bl_43 br_43 wl_39 vdd gnd cell_6t
Xbit_r40_c43 bl_43 br_43 wl_40 vdd gnd cell_6t
Xbit_r41_c43 bl_43 br_43 wl_41 vdd gnd cell_6t
Xbit_r42_c43 bl_43 br_43 wl_42 vdd gnd cell_6t
Xbit_r43_c43 bl_43 br_43 wl_43 vdd gnd cell_6t
Xbit_r44_c43 bl_43 br_43 wl_44 vdd gnd cell_6t
Xbit_r45_c43 bl_43 br_43 wl_45 vdd gnd cell_6t
Xbit_r46_c43 bl_43 br_43 wl_46 vdd gnd cell_6t
Xbit_r47_c43 bl_43 br_43 wl_47 vdd gnd cell_6t
Xbit_r48_c43 bl_43 br_43 wl_48 vdd gnd cell_6t
Xbit_r49_c43 bl_43 br_43 wl_49 vdd gnd cell_6t
Xbit_r50_c43 bl_43 br_43 wl_50 vdd gnd cell_6t
Xbit_r51_c43 bl_43 br_43 wl_51 vdd gnd cell_6t
Xbit_r52_c43 bl_43 br_43 wl_52 vdd gnd cell_6t
Xbit_r53_c43 bl_43 br_43 wl_53 vdd gnd cell_6t
Xbit_r54_c43 bl_43 br_43 wl_54 vdd gnd cell_6t
Xbit_r55_c43 bl_43 br_43 wl_55 vdd gnd cell_6t
Xbit_r56_c43 bl_43 br_43 wl_56 vdd gnd cell_6t
Xbit_r57_c43 bl_43 br_43 wl_57 vdd gnd cell_6t
Xbit_r58_c43 bl_43 br_43 wl_58 vdd gnd cell_6t
Xbit_r59_c43 bl_43 br_43 wl_59 vdd gnd cell_6t
Xbit_r60_c43 bl_43 br_43 wl_60 vdd gnd cell_6t
Xbit_r61_c43 bl_43 br_43 wl_61 vdd gnd cell_6t
Xbit_r62_c43 bl_43 br_43 wl_62 vdd gnd cell_6t
Xbit_r63_c43 bl_43 br_43 wl_63 vdd gnd cell_6t
Xbit_r64_c43 bl_43 br_43 wl_64 vdd gnd cell_6t
Xbit_r65_c43 bl_43 br_43 wl_65 vdd gnd cell_6t
Xbit_r66_c43 bl_43 br_43 wl_66 vdd gnd cell_6t
Xbit_r67_c43 bl_43 br_43 wl_67 vdd gnd cell_6t
Xbit_r68_c43 bl_43 br_43 wl_68 vdd gnd cell_6t
Xbit_r69_c43 bl_43 br_43 wl_69 vdd gnd cell_6t
Xbit_r70_c43 bl_43 br_43 wl_70 vdd gnd cell_6t
Xbit_r71_c43 bl_43 br_43 wl_71 vdd gnd cell_6t
Xbit_r72_c43 bl_43 br_43 wl_72 vdd gnd cell_6t
Xbit_r73_c43 bl_43 br_43 wl_73 vdd gnd cell_6t
Xbit_r74_c43 bl_43 br_43 wl_74 vdd gnd cell_6t
Xbit_r75_c43 bl_43 br_43 wl_75 vdd gnd cell_6t
Xbit_r76_c43 bl_43 br_43 wl_76 vdd gnd cell_6t
Xbit_r77_c43 bl_43 br_43 wl_77 vdd gnd cell_6t
Xbit_r78_c43 bl_43 br_43 wl_78 vdd gnd cell_6t
Xbit_r79_c43 bl_43 br_43 wl_79 vdd gnd cell_6t
Xbit_r80_c43 bl_43 br_43 wl_80 vdd gnd cell_6t
Xbit_r81_c43 bl_43 br_43 wl_81 vdd gnd cell_6t
Xbit_r82_c43 bl_43 br_43 wl_82 vdd gnd cell_6t
Xbit_r83_c43 bl_43 br_43 wl_83 vdd gnd cell_6t
Xbit_r84_c43 bl_43 br_43 wl_84 vdd gnd cell_6t
Xbit_r85_c43 bl_43 br_43 wl_85 vdd gnd cell_6t
Xbit_r86_c43 bl_43 br_43 wl_86 vdd gnd cell_6t
Xbit_r87_c43 bl_43 br_43 wl_87 vdd gnd cell_6t
Xbit_r88_c43 bl_43 br_43 wl_88 vdd gnd cell_6t
Xbit_r89_c43 bl_43 br_43 wl_89 vdd gnd cell_6t
Xbit_r90_c43 bl_43 br_43 wl_90 vdd gnd cell_6t
Xbit_r91_c43 bl_43 br_43 wl_91 vdd gnd cell_6t
Xbit_r92_c43 bl_43 br_43 wl_92 vdd gnd cell_6t
Xbit_r93_c43 bl_43 br_43 wl_93 vdd gnd cell_6t
Xbit_r94_c43 bl_43 br_43 wl_94 vdd gnd cell_6t
Xbit_r95_c43 bl_43 br_43 wl_95 vdd gnd cell_6t
Xbit_r96_c43 bl_43 br_43 wl_96 vdd gnd cell_6t
Xbit_r97_c43 bl_43 br_43 wl_97 vdd gnd cell_6t
Xbit_r98_c43 bl_43 br_43 wl_98 vdd gnd cell_6t
Xbit_r99_c43 bl_43 br_43 wl_99 vdd gnd cell_6t
Xbit_r100_c43 bl_43 br_43 wl_100 vdd gnd cell_6t
Xbit_r101_c43 bl_43 br_43 wl_101 vdd gnd cell_6t
Xbit_r102_c43 bl_43 br_43 wl_102 vdd gnd cell_6t
Xbit_r103_c43 bl_43 br_43 wl_103 vdd gnd cell_6t
Xbit_r104_c43 bl_43 br_43 wl_104 vdd gnd cell_6t
Xbit_r105_c43 bl_43 br_43 wl_105 vdd gnd cell_6t
Xbit_r106_c43 bl_43 br_43 wl_106 vdd gnd cell_6t
Xbit_r107_c43 bl_43 br_43 wl_107 vdd gnd cell_6t
Xbit_r108_c43 bl_43 br_43 wl_108 vdd gnd cell_6t
Xbit_r109_c43 bl_43 br_43 wl_109 vdd gnd cell_6t
Xbit_r110_c43 bl_43 br_43 wl_110 vdd gnd cell_6t
Xbit_r111_c43 bl_43 br_43 wl_111 vdd gnd cell_6t
Xbit_r112_c43 bl_43 br_43 wl_112 vdd gnd cell_6t
Xbit_r113_c43 bl_43 br_43 wl_113 vdd gnd cell_6t
Xbit_r114_c43 bl_43 br_43 wl_114 vdd gnd cell_6t
Xbit_r115_c43 bl_43 br_43 wl_115 vdd gnd cell_6t
Xbit_r116_c43 bl_43 br_43 wl_116 vdd gnd cell_6t
Xbit_r117_c43 bl_43 br_43 wl_117 vdd gnd cell_6t
Xbit_r118_c43 bl_43 br_43 wl_118 vdd gnd cell_6t
Xbit_r119_c43 bl_43 br_43 wl_119 vdd gnd cell_6t
Xbit_r120_c43 bl_43 br_43 wl_120 vdd gnd cell_6t
Xbit_r121_c43 bl_43 br_43 wl_121 vdd gnd cell_6t
Xbit_r122_c43 bl_43 br_43 wl_122 vdd gnd cell_6t
Xbit_r123_c43 bl_43 br_43 wl_123 vdd gnd cell_6t
Xbit_r124_c43 bl_43 br_43 wl_124 vdd gnd cell_6t
Xbit_r125_c43 bl_43 br_43 wl_125 vdd gnd cell_6t
Xbit_r126_c43 bl_43 br_43 wl_126 vdd gnd cell_6t
Xbit_r127_c43 bl_43 br_43 wl_127 vdd gnd cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd cell_6t
Xbit_r1_c44 bl_44 br_44 wl_1 vdd gnd cell_6t
Xbit_r2_c44 bl_44 br_44 wl_2 vdd gnd cell_6t
Xbit_r3_c44 bl_44 br_44 wl_3 vdd gnd cell_6t
Xbit_r4_c44 bl_44 br_44 wl_4 vdd gnd cell_6t
Xbit_r5_c44 bl_44 br_44 wl_5 vdd gnd cell_6t
Xbit_r6_c44 bl_44 br_44 wl_6 vdd gnd cell_6t
Xbit_r7_c44 bl_44 br_44 wl_7 vdd gnd cell_6t
Xbit_r8_c44 bl_44 br_44 wl_8 vdd gnd cell_6t
Xbit_r9_c44 bl_44 br_44 wl_9 vdd gnd cell_6t
Xbit_r10_c44 bl_44 br_44 wl_10 vdd gnd cell_6t
Xbit_r11_c44 bl_44 br_44 wl_11 vdd gnd cell_6t
Xbit_r12_c44 bl_44 br_44 wl_12 vdd gnd cell_6t
Xbit_r13_c44 bl_44 br_44 wl_13 vdd gnd cell_6t
Xbit_r14_c44 bl_44 br_44 wl_14 vdd gnd cell_6t
Xbit_r15_c44 bl_44 br_44 wl_15 vdd gnd cell_6t
Xbit_r16_c44 bl_44 br_44 wl_16 vdd gnd cell_6t
Xbit_r17_c44 bl_44 br_44 wl_17 vdd gnd cell_6t
Xbit_r18_c44 bl_44 br_44 wl_18 vdd gnd cell_6t
Xbit_r19_c44 bl_44 br_44 wl_19 vdd gnd cell_6t
Xbit_r20_c44 bl_44 br_44 wl_20 vdd gnd cell_6t
Xbit_r21_c44 bl_44 br_44 wl_21 vdd gnd cell_6t
Xbit_r22_c44 bl_44 br_44 wl_22 vdd gnd cell_6t
Xbit_r23_c44 bl_44 br_44 wl_23 vdd gnd cell_6t
Xbit_r24_c44 bl_44 br_44 wl_24 vdd gnd cell_6t
Xbit_r25_c44 bl_44 br_44 wl_25 vdd gnd cell_6t
Xbit_r26_c44 bl_44 br_44 wl_26 vdd gnd cell_6t
Xbit_r27_c44 bl_44 br_44 wl_27 vdd gnd cell_6t
Xbit_r28_c44 bl_44 br_44 wl_28 vdd gnd cell_6t
Xbit_r29_c44 bl_44 br_44 wl_29 vdd gnd cell_6t
Xbit_r30_c44 bl_44 br_44 wl_30 vdd gnd cell_6t
Xbit_r31_c44 bl_44 br_44 wl_31 vdd gnd cell_6t
Xbit_r32_c44 bl_44 br_44 wl_32 vdd gnd cell_6t
Xbit_r33_c44 bl_44 br_44 wl_33 vdd gnd cell_6t
Xbit_r34_c44 bl_44 br_44 wl_34 vdd gnd cell_6t
Xbit_r35_c44 bl_44 br_44 wl_35 vdd gnd cell_6t
Xbit_r36_c44 bl_44 br_44 wl_36 vdd gnd cell_6t
Xbit_r37_c44 bl_44 br_44 wl_37 vdd gnd cell_6t
Xbit_r38_c44 bl_44 br_44 wl_38 vdd gnd cell_6t
Xbit_r39_c44 bl_44 br_44 wl_39 vdd gnd cell_6t
Xbit_r40_c44 bl_44 br_44 wl_40 vdd gnd cell_6t
Xbit_r41_c44 bl_44 br_44 wl_41 vdd gnd cell_6t
Xbit_r42_c44 bl_44 br_44 wl_42 vdd gnd cell_6t
Xbit_r43_c44 bl_44 br_44 wl_43 vdd gnd cell_6t
Xbit_r44_c44 bl_44 br_44 wl_44 vdd gnd cell_6t
Xbit_r45_c44 bl_44 br_44 wl_45 vdd gnd cell_6t
Xbit_r46_c44 bl_44 br_44 wl_46 vdd gnd cell_6t
Xbit_r47_c44 bl_44 br_44 wl_47 vdd gnd cell_6t
Xbit_r48_c44 bl_44 br_44 wl_48 vdd gnd cell_6t
Xbit_r49_c44 bl_44 br_44 wl_49 vdd gnd cell_6t
Xbit_r50_c44 bl_44 br_44 wl_50 vdd gnd cell_6t
Xbit_r51_c44 bl_44 br_44 wl_51 vdd gnd cell_6t
Xbit_r52_c44 bl_44 br_44 wl_52 vdd gnd cell_6t
Xbit_r53_c44 bl_44 br_44 wl_53 vdd gnd cell_6t
Xbit_r54_c44 bl_44 br_44 wl_54 vdd gnd cell_6t
Xbit_r55_c44 bl_44 br_44 wl_55 vdd gnd cell_6t
Xbit_r56_c44 bl_44 br_44 wl_56 vdd gnd cell_6t
Xbit_r57_c44 bl_44 br_44 wl_57 vdd gnd cell_6t
Xbit_r58_c44 bl_44 br_44 wl_58 vdd gnd cell_6t
Xbit_r59_c44 bl_44 br_44 wl_59 vdd gnd cell_6t
Xbit_r60_c44 bl_44 br_44 wl_60 vdd gnd cell_6t
Xbit_r61_c44 bl_44 br_44 wl_61 vdd gnd cell_6t
Xbit_r62_c44 bl_44 br_44 wl_62 vdd gnd cell_6t
Xbit_r63_c44 bl_44 br_44 wl_63 vdd gnd cell_6t
Xbit_r64_c44 bl_44 br_44 wl_64 vdd gnd cell_6t
Xbit_r65_c44 bl_44 br_44 wl_65 vdd gnd cell_6t
Xbit_r66_c44 bl_44 br_44 wl_66 vdd gnd cell_6t
Xbit_r67_c44 bl_44 br_44 wl_67 vdd gnd cell_6t
Xbit_r68_c44 bl_44 br_44 wl_68 vdd gnd cell_6t
Xbit_r69_c44 bl_44 br_44 wl_69 vdd gnd cell_6t
Xbit_r70_c44 bl_44 br_44 wl_70 vdd gnd cell_6t
Xbit_r71_c44 bl_44 br_44 wl_71 vdd gnd cell_6t
Xbit_r72_c44 bl_44 br_44 wl_72 vdd gnd cell_6t
Xbit_r73_c44 bl_44 br_44 wl_73 vdd gnd cell_6t
Xbit_r74_c44 bl_44 br_44 wl_74 vdd gnd cell_6t
Xbit_r75_c44 bl_44 br_44 wl_75 vdd gnd cell_6t
Xbit_r76_c44 bl_44 br_44 wl_76 vdd gnd cell_6t
Xbit_r77_c44 bl_44 br_44 wl_77 vdd gnd cell_6t
Xbit_r78_c44 bl_44 br_44 wl_78 vdd gnd cell_6t
Xbit_r79_c44 bl_44 br_44 wl_79 vdd gnd cell_6t
Xbit_r80_c44 bl_44 br_44 wl_80 vdd gnd cell_6t
Xbit_r81_c44 bl_44 br_44 wl_81 vdd gnd cell_6t
Xbit_r82_c44 bl_44 br_44 wl_82 vdd gnd cell_6t
Xbit_r83_c44 bl_44 br_44 wl_83 vdd gnd cell_6t
Xbit_r84_c44 bl_44 br_44 wl_84 vdd gnd cell_6t
Xbit_r85_c44 bl_44 br_44 wl_85 vdd gnd cell_6t
Xbit_r86_c44 bl_44 br_44 wl_86 vdd gnd cell_6t
Xbit_r87_c44 bl_44 br_44 wl_87 vdd gnd cell_6t
Xbit_r88_c44 bl_44 br_44 wl_88 vdd gnd cell_6t
Xbit_r89_c44 bl_44 br_44 wl_89 vdd gnd cell_6t
Xbit_r90_c44 bl_44 br_44 wl_90 vdd gnd cell_6t
Xbit_r91_c44 bl_44 br_44 wl_91 vdd gnd cell_6t
Xbit_r92_c44 bl_44 br_44 wl_92 vdd gnd cell_6t
Xbit_r93_c44 bl_44 br_44 wl_93 vdd gnd cell_6t
Xbit_r94_c44 bl_44 br_44 wl_94 vdd gnd cell_6t
Xbit_r95_c44 bl_44 br_44 wl_95 vdd gnd cell_6t
Xbit_r96_c44 bl_44 br_44 wl_96 vdd gnd cell_6t
Xbit_r97_c44 bl_44 br_44 wl_97 vdd gnd cell_6t
Xbit_r98_c44 bl_44 br_44 wl_98 vdd gnd cell_6t
Xbit_r99_c44 bl_44 br_44 wl_99 vdd gnd cell_6t
Xbit_r100_c44 bl_44 br_44 wl_100 vdd gnd cell_6t
Xbit_r101_c44 bl_44 br_44 wl_101 vdd gnd cell_6t
Xbit_r102_c44 bl_44 br_44 wl_102 vdd gnd cell_6t
Xbit_r103_c44 bl_44 br_44 wl_103 vdd gnd cell_6t
Xbit_r104_c44 bl_44 br_44 wl_104 vdd gnd cell_6t
Xbit_r105_c44 bl_44 br_44 wl_105 vdd gnd cell_6t
Xbit_r106_c44 bl_44 br_44 wl_106 vdd gnd cell_6t
Xbit_r107_c44 bl_44 br_44 wl_107 vdd gnd cell_6t
Xbit_r108_c44 bl_44 br_44 wl_108 vdd gnd cell_6t
Xbit_r109_c44 bl_44 br_44 wl_109 vdd gnd cell_6t
Xbit_r110_c44 bl_44 br_44 wl_110 vdd gnd cell_6t
Xbit_r111_c44 bl_44 br_44 wl_111 vdd gnd cell_6t
Xbit_r112_c44 bl_44 br_44 wl_112 vdd gnd cell_6t
Xbit_r113_c44 bl_44 br_44 wl_113 vdd gnd cell_6t
Xbit_r114_c44 bl_44 br_44 wl_114 vdd gnd cell_6t
Xbit_r115_c44 bl_44 br_44 wl_115 vdd gnd cell_6t
Xbit_r116_c44 bl_44 br_44 wl_116 vdd gnd cell_6t
Xbit_r117_c44 bl_44 br_44 wl_117 vdd gnd cell_6t
Xbit_r118_c44 bl_44 br_44 wl_118 vdd gnd cell_6t
Xbit_r119_c44 bl_44 br_44 wl_119 vdd gnd cell_6t
Xbit_r120_c44 bl_44 br_44 wl_120 vdd gnd cell_6t
Xbit_r121_c44 bl_44 br_44 wl_121 vdd gnd cell_6t
Xbit_r122_c44 bl_44 br_44 wl_122 vdd gnd cell_6t
Xbit_r123_c44 bl_44 br_44 wl_123 vdd gnd cell_6t
Xbit_r124_c44 bl_44 br_44 wl_124 vdd gnd cell_6t
Xbit_r125_c44 bl_44 br_44 wl_125 vdd gnd cell_6t
Xbit_r126_c44 bl_44 br_44 wl_126 vdd gnd cell_6t
Xbit_r127_c44 bl_44 br_44 wl_127 vdd gnd cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd cell_6t
Xbit_r1_c45 bl_45 br_45 wl_1 vdd gnd cell_6t
Xbit_r2_c45 bl_45 br_45 wl_2 vdd gnd cell_6t
Xbit_r3_c45 bl_45 br_45 wl_3 vdd gnd cell_6t
Xbit_r4_c45 bl_45 br_45 wl_4 vdd gnd cell_6t
Xbit_r5_c45 bl_45 br_45 wl_5 vdd gnd cell_6t
Xbit_r6_c45 bl_45 br_45 wl_6 vdd gnd cell_6t
Xbit_r7_c45 bl_45 br_45 wl_7 vdd gnd cell_6t
Xbit_r8_c45 bl_45 br_45 wl_8 vdd gnd cell_6t
Xbit_r9_c45 bl_45 br_45 wl_9 vdd gnd cell_6t
Xbit_r10_c45 bl_45 br_45 wl_10 vdd gnd cell_6t
Xbit_r11_c45 bl_45 br_45 wl_11 vdd gnd cell_6t
Xbit_r12_c45 bl_45 br_45 wl_12 vdd gnd cell_6t
Xbit_r13_c45 bl_45 br_45 wl_13 vdd gnd cell_6t
Xbit_r14_c45 bl_45 br_45 wl_14 vdd gnd cell_6t
Xbit_r15_c45 bl_45 br_45 wl_15 vdd gnd cell_6t
Xbit_r16_c45 bl_45 br_45 wl_16 vdd gnd cell_6t
Xbit_r17_c45 bl_45 br_45 wl_17 vdd gnd cell_6t
Xbit_r18_c45 bl_45 br_45 wl_18 vdd gnd cell_6t
Xbit_r19_c45 bl_45 br_45 wl_19 vdd gnd cell_6t
Xbit_r20_c45 bl_45 br_45 wl_20 vdd gnd cell_6t
Xbit_r21_c45 bl_45 br_45 wl_21 vdd gnd cell_6t
Xbit_r22_c45 bl_45 br_45 wl_22 vdd gnd cell_6t
Xbit_r23_c45 bl_45 br_45 wl_23 vdd gnd cell_6t
Xbit_r24_c45 bl_45 br_45 wl_24 vdd gnd cell_6t
Xbit_r25_c45 bl_45 br_45 wl_25 vdd gnd cell_6t
Xbit_r26_c45 bl_45 br_45 wl_26 vdd gnd cell_6t
Xbit_r27_c45 bl_45 br_45 wl_27 vdd gnd cell_6t
Xbit_r28_c45 bl_45 br_45 wl_28 vdd gnd cell_6t
Xbit_r29_c45 bl_45 br_45 wl_29 vdd gnd cell_6t
Xbit_r30_c45 bl_45 br_45 wl_30 vdd gnd cell_6t
Xbit_r31_c45 bl_45 br_45 wl_31 vdd gnd cell_6t
Xbit_r32_c45 bl_45 br_45 wl_32 vdd gnd cell_6t
Xbit_r33_c45 bl_45 br_45 wl_33 vdd gnd cell_6t
Xbit_r34_c45 bl_45 br_45 wl_34 vdd gnd cell_6t
Xbit_r35_c45 bl_45 br_45 wl_35 vdd gnd cell_6t
Xbit_r36_c45 bl_45 br_45 wl_36 vdd gnd cell_6t
Xbit_r37_c45 bl_45 br_45 wl_37 vdd gnd cell_6t
Xbit_r38_c45 bl_45 br_45 wl_38 vdd gnd cell_6t
Xbit_r39_c45 bl_45 br_45 wl_39 vdd gnd cell_6t
Xbit_r40_c45 bl_45 br_45 wl_40 vdd gnd cell_6t
Xbit_r41_c45 bl_45 br_45 wl_41 vdd gnd cell_6t
Xbit_r42_c45 bl_45 br_45 wl_42 vdd gnd cell_6t
Xbit_r43_c45 bl_45 br_45 wl_43 vdd gnd cell_6t
Xbit_r44_c45 bl_45 br_45 wl_44 vdd gnd cell_6t
Xbit_r45_c45 bl_45 br_45 wl_45 vdd gnd cell_6t
Xbit_r46_c45 bl_45 br_45 wl_46 vdd gnd cell_6t
Xbit_r47_c45 bl_45 br_45 wl_47 vdd gnd cell_6t
Xbit_r48_c45 bl_45 br_45 wl_48 vdd gnd cell_6t
Xbit_r49_c45 bl_45 br_45 wl_49 vdd gnd cell_6t
Xbit_r50_c45 bl_45 br_45 wl_50 vdd gnd cell_6t
Xbit_r51_c45 bl_45 br_45 wl_51 vdd gnd cell_6t
Xbit_r52_c45 bl_45 br_45 wl_52 vdd gnd cell_6t
Xbit_r53_c45 bl_45 br_45 wl_53 vdd gnd cell_6t
Xbit_r54_c45 bl_45 br_45 wl_54 vdd gnd cell_6t
Xbit_r55_c45 bl_45 br_45 wl_55 vdd gnd cell_6t
Xbit_r56_c45 bl_45 br_45 wl_56 vdd gnd cell_6t
Xbit_r57_c45 bl_45 br_45 wl_57 vdd gnd cell_6t
Xbit_r58_c45 bl_45 br_45 wl_58 vdd gnd cell_6t
Xbit_r59_c45 bl_45 br_45 wl_59 vdd gnd cell_6t
Xbit_r60_c45 bl_45 br_45 wl_60 vdd gnd cell_6t
Xbit_r61_c45 bl_45 br_45 wl_61 vdd gnd cell_6t
Xbit_r62_c45 bl_45 br_45 wl_62 vdd gnd cell_6t
Xbit_r63_c45 bl_45 br_45 wl_63 vdd gnd cell_6t
Xbit_r64_c45 bl_45 br_45 wl_64 vdd gnd cell_6t
Xbit_r65_c45 bl_45 br_45 wl_65 vdd gnd cell_6t
Xbit_r66_c45 bl_45 br_45 wl_66 vdd gnd cell_6t
Xbit_r67_c45 bl_45 br_45 wl_67 vdd gnd cell_6t
Xbit_r68_c45 bl_45 br_45 wl_68 vdd gnd cell_6t
Xbit_r69_c45 bl_45 br_45 wl_69 vdd gnd cell_6t
Xbit_r70_c45 bl_45 br_45 wl_70 vdd gnd cell_6t
Xbit_r71_c45 bl_45 br_45 wl_71 vdd gnd cell_6t
Xbit_r72_c45 bl_45 br_45 wl_72 vdd gnd cell_6t
Xbit_r73_c45 bl_45 br_45 wl_73 vdd gnd cell_6t
Xbit_r74_c45 bl_45 br_45 wl_74 vdd gnd cell_6t
Xbit_r75_c45 bl_45 br_45 wl_75 vdd gnd cell_6t
Xbit_r76_c45 bl_45 br_45 wl_76 vdd gnd cell_6t
Xbit_r77_c45 bl_45 br_45 wl_77 vdd gnd cell_6t
Xbit_r78_c45 bl_45 br_45 wl_78 vdd gnd cell_6t
Xbit_r79_c45 bl_45 br_45 wl_79 vdd gnd cell_6t
Xbit_r80_c45 bl_45 br_45 wl_80 vdd gnd cell_6t
Xbit_r81_c45 bl_45 br_45 wl_81 vdd gnd cell_6t
Xbit_r82_c45 bl_45 br_45 wl_82 vdd gnd cell_6t
Xbit_r83_c45 bl_45 br_45 wl_83 vdd gnd cell_6t
Xbit_r84_c45 bl_45 br_45 wl_84 vdd gnd cell_6t
Xbit_r85_c45 bl_45 br_45 wl_85 vdd gnd cell_6t
Xbit_r86_c45 bl_45 br_45 wl_86 vdd gnd cell_6t
Xbit_r87_c45 bl_45 br_45 wl_87 vdd gnd cell_6t
Xbit_r88_c45 bl_45 br_45 wl_88 vdd gnd cell_6t
Xbit_r89_c45 bl_45 br_45 wl_89 vdd gnd cell_6t
Xbit_r90_c45 bl_45 br_45 wl_90 vdd gnd cell_6t
Xbit_r91_c45 bl_45 br_45 wl_91 vdd gnd cell_6t
Xbit_r92_c45 bl_45 br_45 wl_92 vdd gnd cell_6t
Xbit_r93_c45 bl_45 br_45 wl_93 vdd gnd cell_6t
Xbit_r94_c45 bl_45 br_45 wl_94 vdd gnd cell_6t
Xbit_r95_c45 bl_45 br_45 wl_95 vdd gnd cell_6t
Xbit_r96_c45 bl_45 br_45 wl_96 vdd gnd cell_6t
Xbit_r97_c45 bl_45 br_45 wl_97 vdd gnd cell_6t
Xbit_r98_c45 bl_45 br_45 wl_98 vdd gnd cell_6t
Xbit_r99_c45 bl_45 br_45 wl_99 vdd gnd cell_6t
Xbit_r100_c45 bl_45 br_45 wl_100 vdd gnd cell_6t
Xbit_r101_c45 bl_45 br_45 wl_101 vdd gnd cell_6t
Xbit_r102_c45 bl_45 br_45 wl_102 vdd gnd cell_6t
Xbit_r103_c45 bl_45 br_45 wl_103 vdd gnd cell_6t
Xbit_r104_c45 bl_45 br_45 wl_104 vdd gnd cell_6t
Xbit_r105_c45 bl_45 br_45 wl_105 vdd gnd cell_6t
Xbit_r106_c45 bl_45 br_45 wl_106 vdd gnd cell_6t
Xbit_r107_c45 bl_45 br_45 wl_107 vdd gnd cell_6t
Xbit_r108_c45 bl_45 br_45 wl_108 vdd gnd cell_6t
Xbit_r109_c45 bl_45 br_45 wl_109 vdd gnd cell_6t
Xbit_r110_c45 bl_45 br_45 wl_110 vdd gnd cell_6t
Xbit_r111_c45 bl_45 br_45 wl_111 vdd gnd cell_6t
Xbit_r112_c45 bl_45 br_45 wl_112 vdd gnd cell_6t
Xbit_r113_c45 bl_45 br_45 wl_113 vdd gnd cell_6t
Xbit_r114_c45 bl_45 br_45 wl_114 vdd gnd cell_6t
Xbit_r115_c45 bl_45 br_45 wl_115 vdd gnd cell_6t
Xbit_r116_c45 bl_45 br_45 wl_116 vdd gnd cell_6t
Xbit_r117_c45 bl_45 br_45 wl_117 vdd gnd cell_6t
Xbit_r118_c45 bl_45 br_45 wl_118 vdd gnd cell_6t
Xbit_r119_c45 bl_45 br_45 wl_119 vdd gnd cell_6t
Xbit_r120_c45 bl_45 br_45 wl_120 vdd gnd cell_6t
Xbit_r121_c45 bl_45 br_45 wl_121 vdd gnd cell_6t
Xbit_r122_c45 bl_45 br_45 wl_122 vdd gnd cell_6t
Xbit_r123_c45 bl_45 br_45 wl_123 vdd gnd cell_6t
Xbit_r124_c45 bl_45 br_45 wl_124 vdd gnd cell_6t
Xbit_r125_c45 bl_45 br_45 wl_125 vdd gnd cell_6t
Xbit_r126_c45 bl_45 br_45 wl_126 vdd gnd cell_6t
Xbit_r127_c45 bl_45 br_45 wl_127 vdd gnd cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd cell_6t
Xbit_r1_c46 bl_46 br_46 wl_1 vdd gnd cell_6t
Xbit_r2_c46 bl_46 br_46 wl_2 vdd gnd cell_6t
Xbit_r3_c46 bl_46 br_46 wl_3 vdd gnd cell_6t
Xbit_r4_c46 bl_46 br_46 wl_4 vdd gnd cell_6t
Xbit_r5_c46 bl_46 br_46 wl_5 vdd gnd cell_6t
Xbit_r6_c46 bl_46 br_46 wl_6 vdd gnd cell_6t
Xbit_r7_c46 bl_46 br_46 wl_7 vdd gnd cell_6t
Xbit_r8_c46 bl_46 br_46 wl_8 vdd gnd cell_6t
Xbit_r9_c46 bl_46 br_46 wl_9 vdd gnd cell_6t
Xbit_r10_c46 bl_46 br_46 wl_10 vdd gnd cell_6t
Xbit_r11_c46 bl_46 br_46 wl_11 vdd gnd cell_6t
Xbit_r12_c46 bl_46 br_46 wl_12 vdd gnd cell_6t
Xbit_r13_c46 bl_46 br_46 wl_13 vdd gnd cell_6t
Xbit_r14_c46 bl_46 br_46 wl_14 vdd gnd cell_6t
Xbit_r15_c46 bl_46 br_46 wl_15 vdd gnd cell_6t
Xbit_r16_c46 bl_46 br_46 wl_16 vdd gnd cell_6t
Xbit_r17_c46 bl_46 br_46 wl_17 vdd gnd cell_6t
Xbit_r18_c46 bl_46 br_46 wl_18 vdd gnd cell_6t
Xbit_r19_c46 bl_46 br_46 wl_19 vdd gnd cell_6t
Xbit_r20_c46 bl_46 br_46 wl_20 vdd gnd cell_6t
Xbit_r21_c46 bl_46 br_46 wl_21 vdd gnd cell_6t
Xbit_r22_c46 bl_46 br_46 wl_22 vdd gnd cell_6t
Xbit_r23_c46 bl_46 br_46 wl_23 vdd gnd cell_6t
Xbit_r24_c46 bl_46 br_46 wl_24 vdd gnd cell_6t
Xbit_r25_c46 bl_46 br_46 wl_25 vdd gnd cell_6t
Xbit_r26_c46 bl_46 br_46 wl_26 vdd gnd cell_6t
Xbit_r27_c46 bl_46 br_46 wl_27 vdd gnd cell_6t
Xbit_r28_c46 bl_46 br_46 wl_28 vdd gnd cell_6t
Xbit_r29_c46 bl_46 br_46 wl_29 vdd gnd cell_6t
Xbit_r30_c46 bl_46 br_46 wl_30 vdd gnd cell_6t
Xbit_r31_c46 bl_46 br_46 wl_31 vdd gnd cell_6t
Xbit_r32_c46 bl_46 br_46 wl_32 vdd gnd cell_6t
Xbit_r33_c46 bl_46 br_46 wl_33 vdd gnd cell_6t
Xbit_r34_c46 bl_46 br_46 wl_34 vdd gnd cell_6t
Xbit_r35_c46 bl_46 br_46 wl_35 vdd gnd cell_6t
Xbit_r36_c46 bl_46 br_46 wl_36 vdd gnd cell_6t
Xbit_r37_c46 bl_46 br_46 wl_37 vdd gnd cell_6t
Xbit_r38_c46 bl_46 br_46 wl_38 vdd gnd cell_6t
Xbit_r39_c46 bl_46 br_46 wl_39 vdd gnd cell_6t
Xbit_r40_c46 bl_46 br_46 wl_40 vdd gnd cell_6t
Xbit_r41_c46 bl_46 br_46 wl_41 vdd gnd cell_6t
Xbit_r42_c46 bl_46 br_46 wl_42 vdd gnd cell_6t
Xbit_r43_c46 bl_46 br_46 wl_43 vdd gnd cell_6t
Xbit_r44_c46 bl_46 br_46 wl_44 vdd gnd cell_6t
Xbit_r45_c46 bl_46 br_46 wl_45 vdd gnd cell_6t
Xbit_r46_c46 bl_46 br_46 wl_46 vdd gnd cell_6t
Xbit_r47_c46 bl_46 br_46 wl_47 vdd gnd cell_6t
Xbit_r48_c46 bl_46 br_46 wl_48 vdd gnd cell_6t
Xbit_r49_c46 bl_46 br_46 wl_49 vdd gnd cell_6t
Xbit_r50_c46 bl_46 br_46 wl_50 vdd gnd cell_6t
Xbit_r51_c46 bl_46 br_46 wl_51 vdd gnd cell_6t
Xbit_r52_c46 bl_46 br_46 wl_52 vdd gnd cell_6t
Xbit_r53_c46 bl_46 br_46 wl_53 vdd gnd cell_6t
Xbit_r54_c46 bl_46 br_46 wl_54 vdd gnd cell_6t
Xbit_r55_c46 bl_46 br_46 wl_55 vdd gnd cell_6t
Xbit_r56_c46 bl_46 br_46 wl_56 vdd gnd cell_6t
Xbit_r57_c46 bl_46 br_46 wl_57 vdd gnd cell_6t
Xbit_r58_c46 bl_46 br_46 wl_58 vdd gnd cell_6t
Xbit_r59_c46 bl_46 br_46 wl_59 vdd gnd cell_6t
Xbit_r60_c46 bl_46 br_46 wl_60 vdd gnd cell_6t
Xbit_r61_c46 bl_46 br_46 wl_61 vdd gnd cell_6t
Xbit_r62_c46 bl_46 br_46 wl_62 vdd gnd cell_6t
Xbit_r63_c46 bl_46 br_46 wl_63 vdd gnd cell_6t
Xbit_r64_c46 bl_46 br_46 wl_64 vdd gnd cell_6t
Xbit_r65_c46 bl_46 br_46 wl_65 vdd gnd cell_6t
Xbit_r66_c46 bl_46 br_46 wl_66 vdd gnd cell_6t
Xbit_r67_c46 bl_46 br_46 wl_67 vdd gnd cell_6t
Xbit_r68_c46 bl_46 br_46 wl_68 vdd gnd cell_6t
Xbit_r69_c46 bl_46 br_46 wl_69 vdd gnd cell_6t
Xbit_r70_c46 bl_46 br_46 wl_70 vdd gnd cell_6t
Xbit_r71_c46 bl_46 br_46 wl_71 vdd gnd cell_6t
Xbit_r72_c46 bl_46 br_46 wl_72 vdd gnd cell_6t
Xbit_r73_c46 bl_46 br_46 wl_73 vdd gnd cell_6t
Xbit_r74_c46 bl_46 br_46 wl_74 vdd gnd cell_6t
Xbit_r75_c46 bl_46 br_46 wl_75 vdd gnd cell_6t
Xbit_r76_c46 bl_46 br_46 wl_76 vdd gnd cell_6t
Xbit_r77_c46 bl_46 br_46 wl_77 vdd gnd cell_6t
Xbit_r78_c46 bl_46 br_46 wl_78 vdd gnd cell_6t
Xbit_r79_c46 bl_46 br_46 wl_79 vdd gnd cell_6t
Xbit_r80_c46 bl_46 br_46 wl_80 vdd gnd cell_6t
Xbit_r81_c46 bl_46 br_46 wl_81 vdd gnd cell_6t
Xbit_r82_c46 bl_46 br_46 wl_82 vdd gnd cell_6t
Xbit_r83_c46 bl_46 br_46 wl_83 vdd gnd cell_6t
Xbit_r84_c46 bl_46 br_46 wl_84 vdd gnd cell_6t
Xbit_r85_c46 bl_46 br_46 wl_85 vdd gnd cell_6t
Xbit_r86_c46 bl_46 br_46 wl_86 vdd gnd cell_6t
Xbit_r87_c46 bl_46 br_46 wl_87 vdd gnd cell_6t
Xbit_r88_c46 bl_46 br_46 wl_88 vdd gnd cell_6t
Xbit_r89_c46 bl_46 br_46 wl_89 vdd gnd cell_6t
Xbit_r90_c46 bl_46 br_46 wl_90 vdd gnd cell_6t
Xbit_r91_c46 bl_46 br_46 wl_91 vdd gnd cell_6t
Xbit_r92_c46 bl_46 br_46 wl_92 vdd gnd cell_6t
Xbit_r93_c46 bl_46 br_46 wl_93 vdd gnd cell_6t
Xbit_r94_c46 bl_46 br_46 wl_94 vdd gnd cell_6t
Xbit_r95_c46 bl_46 br_46 wl_95 vdd gnd cell_6t
Xbit_r96_c46 bl_46 br_46 wl_96 vdd gnd cell_6t
Xbit_r97_c46 bl_46 br_46 wl_97 vdd gnd cell_6t
Xbit_r98_c46 bl_46 br_46 wl_98 vdd gnd cell_6t
Xbit_r99_c46 bl_46 br_46 wl_99 vdd gnd cell_6t
Xbit_r100_c46 bl_46 br_46 wl_100 vdd gnd cell_6t
Xbit_r101_c46 bl_46 br_46 wl_101 vdd gnd cell_6t
Xbit_r102_c46 bl_46 br_46 wl_102 vdd gnd cell_6t
Xbit_r103_c46 bl_46 br_46 wl_103 vdd gnd cell_6t
Xbit_r104_c46 bl_46 br_46 wl_104 vdd gnd cell_6t
Xbit_r105_c46 bl_46 br_46 wl_105 vdd gnd cell_6t
Xbit_r106_c46 bl_46 br_46 wl_106 vdd gnd cell_6t
Xbit_r107_c46 bl_46 br_46 wl_107 vdd gnd cell_6t
Xbit_r108_c46 bl_46 br_46 wl_108 vdd gnd cell_6t
Xbit_r109_c46 bl_46 br_46 wl_109 vdd gnd cell_6t
Xbit_r110_c46 bl_46 br_46 wl_110 vdd gnd cell_6t
Xbit_r111_c46 bl_46 br_46 wl_111 vdd gnd cell_6t
Xbit_r112_c46 bl_46 br_46 wl_112 vdd gnd cell_6t
Xbit_r113_c46 bl_46 br_46 wl_113 vdd gnd cell_6t
Xbit_r114_c46 bl_46 br_46 wl_114 vdd gnd cell_6t
Xbit_r115_c46 bl_46 br_46 wl_115 vdd gnd cell_6t
Xbit_r116_c46 bl_46 br_46 wl_116 vdd gnd cell_6t
Xbit_r117_c46 bl_46 br_46 wl_117 vdd gnd cell_6t
Xbit_r118_c46 bl_46 br_46 wl_118 vdd gnd cell_6t
Xbit_r119_c46 bl_46 br_46 wl_119 vdd gnd cell_6t
Xbit_r120_c46 bl_46 br_46 wl_120 vdd gnd cell_6t
Xbit_r121_c46 bl_46 br_46 wl_121 vdd gnd cell_6t
Xbit_r122_c46 bl_46 br_46 wl_122 vdd gnd cell_6t
Xbit_r123_c46 bl_46 br_46 wl_123 vdd gnd cell_6t
Xbit_r124_c46 bl_46 br_46 wl_124 vdd gnd cell_6t
Xbit_r125_c46 bl_46 br_46 wl_125 vdd gnd cell_6t
Xbit_r126_c46 bl_46 br_46 wl_126 vdd gnd cell_6t
Xbit_r127_c46 bl_46 br_46 wl_127 vdd gnd cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd cell_6t
Xbit_r1_c47 bl_47 br_47 wl_1 vdd gnd cell_6t
Xbit_r2_c47 bl_47 br_47 wl_2 vdd gnd cell_6t
Xbit_r3_c47 bl_47 br_47 wl_3 vdd gnd cell_6t
Xbit_r4_c47 bl_47 br_47 wl_4 vdd gnd cell_6t
Xbit_r5_c47 bl_47 br_47 wl_5 vdd gnd cell_6t
Xbit_r6_c47 bl_47 br_47 wl_6 vdd gnd cell_6t
Xbit_r7_c47 bl_47 br_47 wl_7 vdd gnd cell_6t
Xbit_r8_c47 bl_47 br_47 wl_8 vdd gnd cell_6t
Xbit_r9_c47 bl_47 br_47 wl_9 vdd gnd cell_6t
Xbit_r10_c47 bl_47 br_47 wl_10 vdd gnd cell_6t
Xbit_r11_c47 bl_47 br_47 wl_11 vdd gnd cell_6t
Xbit_r12_c47 bl_47 br_47 wl_12 vdd gnd cell_6t
Xbit_r13_c47 bl_47 br_47 wl_13 vdd gnd cell_6t
Xbit_r14_c47 bl_47 br_47 wl_14 vdd gnd cell_6t
Xbit_r15_c47 bl_47 br_47 wl_15 vdd gnd cell_6t
Xbit_r16_c47 bl_47 br_47 wl_16 vdd gnd cell_6t
Xbit_r17_c47 bl_47 br_47 wl_17 vdd gnd cell_6t
Xbit_r18_c47 bl_47 br_47 wl_18 vdd gnd cell_6t
Xbit_r19_c47 bl_47 br_47 wl_19 vdd gnd cell_6t
Xbit_r20_c47 bl_47 br_47 wl_20 vdd gnd cell_6t
Xbit_r21_c47 bl_47 br_47 wl_21 vdd gnd cell_6t
Xbit_r22_c47 bl_47 br_47 wl_22 vdd gnd cell_6t
Xbit_r23_c47 bl_47 br_47 wl_23 vdd gnd cell_6t
Xbit_r24_c47 bl_47 br_47 wl_24 vdd gnd cell_6t
Xbit_r25_c47 bl_47 br_47 wl_25 vdd gnd cell_6t
Xbit_r26_c47 bl_47 br_47 wl_26 vdd gnd cell_6t
Xbit_r27_c47 bl_47 br_47 wl_27 vdd gnd cell_6t
Xbit_r28_c47 bl_47 br_47 wl_28 vdd gnd cell_6t
Xbit_r29_c47 bl_47 br_47 wl_29 vdd gnd cell_6t
Xbit_r30_c47 bl_47 br_47 wl_30 vdd gnd cell_6t
Xbit_r31_c47 bl_47 br_47 wl_31 vdd gnd cell_6t
Xbit_r32_c47 bl_47 br_47 wl_32 vdd gnd cell_6t
Xbit_r33_c47 bl_47 br_47 wl_33 vdd gnd cell_6t
Xbit_r34_c47 bl_47 br_47 wl_34 vdd gnd cell_6t
Xbit_r35_c47 bl_47 br_47 wl_35 vdd gnd cell_6t
Xbit_r36_c47 bl_47 br_47 wl_36 vdd gnd cell_6t
Xbit_r37_c47 bl_47 br_47 wl_37 vdd gnd cell_6t
Xbit_r38_c47 bl_47 br_47 wl_38 vdd gnd cell_6t
Xbit_r39_c47 bl_47 br_47 wl_39 vdd gnd cell_6t
Xbit_r40_c47 bl_47 br_47 wl_40 vdd gnd cell_6t
Xbit_r41_c47 bl_47 br_47 wl_41 vdd gnd cell_6t
Xbit_r42_c47 bl_47 br_47 wl_42 vdd gnd cell_6t
Xbit_r43_c47 bl_47 br_47 wl_43 vdd gnd cell_6t
Xbit_r44_c47 bl_47 br_47 wl_44 vdd gnd cell_6t
Xbit_r45_c47 bl_47 br_47 wl_45 vdd gnd cell_6t
Xbit_r46_c47 bl_47 br_47 wl_46 vdd gnd cell_6t
Xbit_r47_c47 bl_47 br_47 wl_47 vdd gnd cell_6t
Xbit_r48_c47 bl_47 br_47 wl_48 vdd gnd cell_6t
Xbit_r49_c47 bl_47 br_47 wl_49 vdd gnd cell_6t
Xbit_r50_c47 bl_47 br_47 wl_50 vdd gnd cell_6t
Xbit_r51_c47 bl_47 br_47 wl_51 vdd gnd cell_6t
Xbit_r52_c47 bl_47 br_47 wl_52 vdd gnd cell_6t
Xbit_r53_c47 bl_47 br_47 wl_53 vdd gnd cell_6t
Xbit_r54_c47 bl_47 br_47 wl_54 vdd gnd cell_6t
Xbit_r55_c47 bl_47 br_47 wl_55 vdd gnd cell_6t
Xbit_r56_c47 bl_47 br_47 wl_56 vdd gnd cell_6t
Xbit_r57_c47 bl_47 br_47 wl_57 vdd gnd cell_6t
Xbit_r58_c47 bl_47 br_47 wl_58 vdd gnd cell_6t
Xbit_r59_c47 bl_47 br_47 wl_59 vdd gnd cell_6t
Xbit_r60_c47 bl_47 br_47 wl_60 vdd gnd cell_6t
Xbit_r61_c47 bl_47 br_47 wl_61 vdd gnd cell_6t
Xbit_r62_c47 bl_47 br_47 wl_62 vdd gnd cell_6t
Xbit_r63_c47 bl_47 br_47 wl_63 vdd gnd cell_6t
Xbit_r64_c47 bl_47 br_47 wl_64 vdd gnd cell_6t
Xbit_r65_c47 bl_47 br_47 wl_65 vdd gnd cell_6t
Xbit_r66_c47 bl_47 br_47 wl_66 vdd gnd cell_6t
Xbit_r67_c47 bl_47 br_47 wl_67 vdd gnd cell_6t
Xbit_r68_c47 bl_47 br_47 wl_68 vdd gnd cell_6t
Xbit_r69_c47 bl_47 br_47 wl_69 vdd gnd cell_6t
Xbit_r70_c47 bl_47 br_47 wl_70 vdd gnd cell_6t
Xbit_r71_c47 bl_47 br_47 wl_71 vdd gnd cell_6t
Xbit_r72_c47 bl_47 br_47 wl_72 vdd gnd cell_6t
Xbit_r73_c47 bl_47 br_47 wl_73 vdd gnd cell_6t
Xbit_r74_c47 bl_47 br_47 wl_74 vdd gnd cell_6t
Xbit_r75_c47 bl_47 br_47 wl_75 vdd gnd cell_6t
Xbit_r76_c47 bl_47 br_47 wl_76 vdd gnd cell_6t
Xbit_r77_c47 bl_47 br_47 wl_77 vdd gnd cell_6t
Xbit_r78_c47 bl_47 br_47 wl_78 vdd gnd cell_6t
Xbit_r79_c47 bl_47 br_47 wl_79 vdd gnd cell_6t
Xbit_r80_c47 bl_47 br_47 wl_80 vdd gnd cell_6t
Xbit_r81_c47 bl_47 br_47 wl_81 vdd gnd cell_6t
Xbit_r82_c47 bl_47 br_47 wl_82 vdd gnd cell_6t
Xbit_r83_c47 bl_47 br_47 wl_83 vdd gnd cell_6t
Xbit_r84_c47 bl_47 br_47 wl_84 vdd gnd cell_6t
Xbit_r85_c47 bl_47 br_47 wl_85 vdd gnd cell_6t
Xbit_r86_c47 bl_47 br_47 wl_86 vdd gnd cell_6t
Xbit_r87_c47 bl_47 br_47 wl_87 vdd gnd cell_6t
Xbit_r88_c47 bl_47 br_47 wl_88 vdd gnd cell_6t
Xbit_r89_c47 bl_47 br_47 wl_89 vdd gnd cell_6t
Xbit_r90_c47 bl_47 br_47 wl_90 vdd gnd cell_6t
Xbit_r91_c47 bl_47 br_47 wl_91 vdd gnd cell_6t
Xbit_r92_c47 bl_47 br_47 wl_92 vdd gnd cell_6t
Xbit_r93_c47 bl_47 br_47 wl_93 vdd gnd cell_6t
Xbit_r94_c47 bl_47 br_47 wl_94 vdd gnd cell_6t
Xbit_r95_c47 bl_47 br_47 wl_95 vdd gnd cell_6t
Xbit_r96_c47 bl_47 br_47 wl_96 vdd gnd cell_6t
Xbit_r97_c47 bl_47 br_47 wl_97 vdd gnd cell_6t
Xbit_r98_c47 bl_47 br_47 wl_98 vdd gnd cell_6t
Xbit_r99_c47 bl_47 br_47 wl_99 vdd gnd cell_6t
Xbit_r100_c47 bl_47 br_47 wl_100 vdd gnd cell_6t
Xbit_r101_c47 bl_47 br_47 wl_101 vdd gnd cell_6t
Xbit_r102_c47 bl_47 br_47 wl_102 vdd gnd cell_6t
Xbit_r103_c47 bl_47 br_47 wl_103 vdd gnd cell_6t
Xbit_r104_c47 bl_47 br_47 wl_104 vdd gnd cell_6t
Xbit_r105_c47 bl_47 br_47 wl_105 vdd gnd cell_6t
Xbit_r106_c47 bl_47 br_47 wl_106 vdd gnd cell_6t
Xbit_r107_c47 bl_47 br_47 wl_107 vdd gnd cell_6t
Xbit_r108_c47 bl_47 br_47 wl_108 vdd gnd cell_6t
Xbit_r109_c47 bl_47 br_47 wl_109 vdd gnd cell_6t
Xbit_r110_c47 bl_47 br_47 wl_110 vdd gnd cell_6t
Xbit_r111_c47 bl_47 br_47 wl_111 vdd gnd cell_6t
Xbit_r112_c47 bl_47 br_47 wl_112 vdd gnd cell_6t
Xbit_r113_c47 bl_47 br_47 wl_113 vdd gnd cell_6t
Xbit_r114_c47 bl_47 br_47 wl_114 vdd gnd cell_6t
Xbit_r115_c47 bl_47 br_47 wl_115 vdd gnd cell_6t
Xbit_r116_c47 bl_47 br_47 wl_116 vdd gnd cell_6t
Xbit_r117_c47 bl_47 br_47 wl_117 vdd gnd cell_6t
Xbit_r118_c47 bl_47 br_47 wl_118 vdd gnd cell_6t
Xbit_r119_c47 bl_47 br_47 wl_119 vdd gnd cell_6t
Xbit_r120_c47 bl_47 br_47 wl_120 vdd gnd cell_6t
Xbit_r121_c47 bl_47 br_47 wl_121 vdd gnd cell_6t
Xbit_r122_c47 bl_47 br_47 wl_122 vdd gnd cell_6t
Xbit_r123_c47 bl_47 br_47 wl_123 vdd gnd cell_6t
Xbit_r124_c47 bl_47 br_47 wl_124 vdd gnd cell_6t
Xbit_r125_c47 bl_47 br_47 wl_125 vdd gnd cell_6t
Xbit_r126_c47 bl_47 br_47 wl_126 vdd gnd cell_6t
Xbit_r127_c47 bl_47 br_47 wl_127 vdd gnd cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd cell_6t
Xbit_r1_c48 bl_48 br_48 wl_1 vdd gnd cell_6t
Xbit_r2_c48 bl_48 br_48 wl_2 vdd gnd cell_6t
Xbit_r3_c48 bl_48 br_48 wl_3 vdd gnd cell_6t
Xbit_r4_c48 bl_48 br_48 wl_4 vdd gnd cell_6t
Xbit_r5_c48 bl_48 br_48 wl_5 vdd gnd cell_6t
Xbit_r6_c48 bl_48 br_48 wl_6 vdd gnd cell_6t
Xbit_r7_c48 bl_48 br_48 wl_7 vdd gnd cell_6t
Xbit_r8_c48 bl_48 br_48 wl_8 vdd gnd cell_6t
Xbit_r9_c48 bl_48 br_48 wl_9 vdd gnd cell_6t
Xbit_r10_c48 bl_48 br_48 wl_10 vdd gnd cell_6t
Xbit_r11_c48 bl_48 br_48 wl_11 vdd gnd cell_6t
Xbit_r12_c48 bl_48 br_48 wl_12 vdd gnd cell_6t
Xbit_r13_c48 bl_48 br_48 wl_13 vdd gnd cell_6t
Xbit_r14_c48 bl_48 br_48 wl_14 vdd gnd cell_6t
Xbit_r15_c48 bl_48 br_48 wl_15 vdd gnd cell_6t
Xbit_r16_c48 bl_48 br_48 wl_16 vdd gnd cell_6t
Xbit_r17_c48 bl_48 br_48 wl_17 vdd gnd cell_6t
Xbit_r18_c48 bl_48 br_48 wl_18 vdd gnd cell_6t
Xbit_r19_c48 bl_48 br_48 wl_19 vdd gnd cell_6t
Xbit_r20_c48 bl_48 br_48 wl_20 vdd gnd cell_6t
Xbit_r21_c48 bl_48 br_48 wl_21 vdd gnd cell_6t
Xbit_r22_c48 bl_48 br_48 wl_22 vdd gnd cell_6t
Xbit_r23_c48 bl_48 br_48 wl_23 vdd gnd cell_6t
Xbit_r24_c48 bl_48 br_48 wl_24 vdd gnd cell_6t
Xbit_r25_c48 bl_48 br_48 wl_25 vdd gnd cell_6t
Xbit_r26_c48 bl_48 br_48 wl_26 vdd gnd cell_6t
Xbit_r27_c48 bl_48 br_48 wl_27 vdd gnd cell_6t
Xbit_r28_c48 bl_48 br_48 wl_28 vdd gnd cell_6t
Xbit_r29_c48 bl_48 br_48 wl_29 vdd gnd cell_6t
Xbit_r30_c48 bl_48 br_48 wl_30 vdd gnd cell_6t
Xbit_r31_c48 bl_48 br_48 wl_31 vdd gnd cell_6t
Xbit_r32_c48 bl_48 br_48 wl_32 vdd gnd cell_6t
Xbit_r33_c48 bl_48 br_48 wl_33 vdd gnd cell_6t
Xbit_r34_c48 bl_48 br_48 wl_34 vdd gnd cell_6t
Xbit_r35_c48 bl_48 br_48 wl_35 vdd gnd cell_6t
Xbit_r36_c48 bl_48 br_48 wl_36 vdd gnd cell_6t
Xbit_r37_c48 bl_48 br_48 wl_37 vdd gnd cell_6t
Xbit_r38_c48 bl_48 br_48 wl_38 vdd gnd cell_6t
Xbit_r39_c48 bl_48 br_48 wl_39 vdd gnd cell_6t
Xbit_r40_c48 bl_48 br_48 wl_40 vdd gnd cell_6t
Xbit_r41_c48 bl_48 br_48 wl_41 vdd gnd cell_6t
Xbit_r42_c48 bl_48 br_48 wl_42 vdd gnd cell_6t
Xbit_r43_c48 bl_48 br_48 wl_43 vdd gnd cell_6t
Xbit_r44_c48 bl_48 br_48 wl_44 vdd gnd cell_6t
Xbit_r45_c48 bl_48 br_48 wl_45 vdd gnd cell_6t
Xbit_r46_c48 bl_48 br_48 wl_46 vdd gnd cell_6t
Xbit_r47_c48 bl_48 br_48 wl_47 vdd gnd cell_6t
Xbit_r48_c48 bl_48 br_48 wl_48 vdd gnd cell_6t
Xbit_r49_c48 bl_48 br_48 wl_49 vdd gnd cell_6t
Xbit_r50_c48 bl_48 br_48 wl_50 vdd gnd cell_6t
Xbit_r51_c48 bl_48 br_48 wl_51 vdd gnd cell_6t
Xbit_r52_c48 bl_48 br_48 wl_52 vdd gnd cell_6t
Xbit_r53_c48 bl_48 br_48 wl_53 vdd gnd cell_6t
Xbit_r54_c48 bl_48 br_48 wl_54 vdd gnd cell_6t
Xbit_r55_c48 bl_48 br_48 wl_55 vdd gnd cell_6t
Xbit_r56_c48 bl_48 br_48 wl_56 vdd gnd cell_6t
Xbit_r57_c48 bl_48 br_48 wl_57 vdd gnd cell_6t
Xbit_r58_c48 bl_48 br_48 wl_58 vdd gnd cell_6t
Xbit_r59_c48 bl_48 br_48 wl_59 vdd gnd cell_6t
Xbit_r60_c48 bl_48 br_48 wl_60 vdd gnd cell_6t
Xbit_r61_c48 bl_48 br_48 wl_61 vdd gnd cell_6t
Xbit_r62_c48 bl_48 br_48 wl_62 vdd gnd cell_6t
Xbit_r63_c48 bl_48 br_48 wl_63 vdd gnd cell_6t
Xbit_r64_c48 bl_48 br_48 wl_64 vdd gnd cell_6t
Xbit_r65_c48 bl_48 br_48 wl_65 vdd gnd cell_6t
Xbit_r66_c48 bl_48 br_48 wl_66 vdd gnd cell_6t
Xbit_r67_c48 bl_48 br_48 wl_67 vdd gnd cell_6t
Xbit_r68_c48 bl_48 br_48 wl_68 vdd gnd cell_6t
Xbit_r69_c48 bl_48 br_48 wl_69 vdd gnd cell_6t
Xbit_r70_c48 bl_48 br_48 wl_70 vdd gnd cell_6t
Xbit_r71_c48 bl_48 br_48 wl_71 vdd gnd cell_6t
Xbit_r72_c48 bl_48 br_48 wl_72 vdd gnd cell_6t
Xbit_r73_c48 bl_48 br_48 wl_73 vdd gnd cell_6t
Xbit_r74_c48 bl_48 br_48 wl_74 vdd gnd cell_6t
Xbit_r75_c48 bl_48 br_48 wl_75 vdd gnd cell_6t
Xbit_r76_c48 bl_48 br_48 wl_76 vdd gnd cell_6t
Xbit_r77_c48 bl_48 br_48 wl_77 vdd gnd cell_6t
Xbit_r78_c48 bl_48 br_48 wl_78 vdd gnd cell_6t
Xbit_r79_c48 bl_48 br_48 wl_79 vdd gnd cell_6t
Xbit_r80_c48 bl_48 br_48 wl_80 vdd gnd cell_6t
Xbit_r81_c48 bl_48 br_48 wl_81 vdd gnd cell_6t
Xbit_r82_c48 bl_48 br_48 wl_82 vdd gnd cell_6t
Xbit_r83_c48 bl_48 br_48 wl_83 vdd gnd cell_6t
Xbit_r84_c48 bl_48 br_48 wl_84 vdd gnd cell_6t
Xbit_r85_c48 bl_48 br_48 wl_85 vdd gnd cell_6t
Xbit_r86_c48 bl_48 br_48 wl_86 vdd gnd cell_6t
Xbit_r87_c48 bl_48 br_48 wl_87 vdd gnd cell_6t
Xbit_r88_c48 bl_48 br_48 wl_88 vdd gnd cell_6t
Xbit_r89_c48 bl_48 br_48 wl_89 vdd gnd cell_6t
Xbit_r90_c48 bl_48 br_48 wl_90 vdd gnd cell_6t
Xbit_r91_c48 bl_48 br_48 wl_91 vdd gnd cell_6t
Xbit_r92_c48 bl_48 br_48 wl_92 vdd gnd cell_6t
Xbit_r93_c48 bl_48 br_48 wl_93 vdd gnd cell_6t
Xbit_r94_c48 bl_48 br_48 wl_94 vdd gnd cell_6t
Xbit_r95_c48 bl_48 br_48 wl_95 vdd gnd cell_6t
Xbit_r96_c48 bl_48 br_48 wl_96 vdd gnd cell_6t
Xbit_r97_c48 bl_48 br_48 wl_97 vdd gnd cell_6t
Xbit_r98_c48 bl_48 br_48 wl_98 vdd gnd cell_6t
Xbit_r99_c48 bl_48 br_48 wl_99 vdd gnd cell_6t
Xbit_r100_c48 bl_48 br_48 wl_100 vdd gnd cell_6t
Xbit_r101_c48 bl_48 br_48 wl_101 vdd gnd cell_6t
Xbit_r102_c48 bl_48 br_48 wl_102 vdd gnd cell_6t
Xbit_r103_c48 bl_48 br_48 wl_103 vdd gnd cell_6t
Xbit_r104_c48 bl_48 br_48 wl_104 vdd gnd cell_6t
Xbit_r105_c48 bl_48 br_48 wl_105 vdd gnd cell_6t
Xbit_r106_c48 bl_48 br_48 wl_106 vdd gnd cell_6t
Xbit_r107_c48 bl_48 br_48 wl_107 vdd gnd cell_6t
Xbit_r108_c48 bl_48 br_48 wl_108 vdd gnd cell_6t
Xbit_r109_c48 bl_48 br_48 wl_109 vdd gnd cell_6t
Xbit_r110_c48 bl_48 br_48 wl_110 vdd gnd cell_6t
Xbit_r111_c48 bl_48 br_48 wl_111 vdd gnd cell_6t
Xbit_r112_c48 bl_48 br_48 wl_112 vdd gnd cell_6t
Xbit_r113_c48 bl_48 br_48 wl_113 vdd gnd cell_6t
Xbit_r114_c48 bl_48 br_48 wl_114 vdd gnd cell_6t
Xbit_r115_c48 bl_48 br_48 wl_115 vdd gnd cell_6t
Xbit_r116_c48 bl_48 br_48 wl_116 vdd gnd cell_6t
Xbit_r117_c48 bl_48 br_48 wl_117 vdd gnd cell_6t
Xbit_r118_c48 bl_48 br_48 wl_118 vdd gnd cell_6t
Xbit_r119_c48 bl_48 br_48 wl_119 vdd gnd cell_6t
Xbit_r120_c48 bl_48 br_48 wl_120 vdd gnd cell_6t
Xbit_r121_c48 bl_48 br_48 wl_121 vdd gnd cell_6t
Xbit_r122_c48 bl_48 br_48 wl_122 vdd gnd cell_6t
Xbit_r123_c48 bl_48 br_48 wl_123 vdd gnd cell_6t
Xbit_r124_c48 bl_48 br_48 wl_124 vdd gnd cell_6t
Xbit_r125_c48 bl_48 br_48 wl_125 vdd gnd cell_6t
Xbit_r126_c48 bl_48 br_48 wl_126 vdd gnd cell_6t
Xbit_r127_c48 bl_48 br_48 wl_127 vdd gnd cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd cell_6t
Xbit_r1_c49 bl_49 br_49 wl_1 vdd gnd cell_6t
Xbit_r2_c49 bl_49 br_49 wl_2 vdd gnd cell_6t
Xbit_r3_c49 bl_49 br_49 wl_3 vdd gnd cell_6t
Xbit_r4_c49 bl_49 br_49 wl_4 vdd gnd cell_6t
Xbit_r5_c49 bl_49 br_49 wl_5 vdd gnd cell_6t
Xbit_r6_c49 bl_49 br_49 wl_6 vdd gnd cell_6t
Xbit_r7_c49 bl_49 br_49 wl_7 vdd gnd cell_6t
Xbit_r8_c49 bl_49 br_49 wl_8 vdd gnd cell_6t
Xbit_r9_c49 bl_49 br_49 wl_9 vdd gnd cell_6t
Xbit_r10_c49 bl_49 br_49 wl_10 vdd gnd cell_6t
Xbit_r11_c49 bl_49 br_49 wl_11 vdd gnd cell_6t
Xbit_r12_c49 bl_49 br_49 wl_12 vdd gnd cell_6t
Xbit_r13_c49 bl_49 br_49 wl_13 vdd gnd cell_6t
Xbit_r14_c49 bl_49 br_49 wl_14 vdd gnd cell_6t
Xbit_r15_c49 bl_49 br_49 wl_15 vdd gnd cell_6t
Xbit_r16_c49 bl_49 br_49 wl_16 vdd gnd cell_6t
Xbit_r17_c49 bl_49 br_49 wl_17 vdd gnd cell_6t
Xbit_r18_c49 bl_49 br_49 wl_18 vdd gnd cell_6t
Xbit_r19_c49 bl_49 br_49 wl_19 vdd gnd cell_6t
Xbit_r20_c49 bl_49 br_49 wl_20 vdd gnd cell_6t
Xbit_r21_c49 bl_49 br_49 wl_21 vdd gnd cell_6t
Xbit_r22_c49 bl_49 br_49 wl_22 vdd gnd cell_6t
Xbit_r23_c49 bl_49 br_49 wl_23 vdd gnd cell_6t
Xbit_r24_c49 bl_49 br_49 wl_24 vdd gnd cell_6t
Xbit_r25_c49 bl_49 br_49 wl_25 vdd gnd cell_6t
Xbit_r26_c49 bl_49 br_49 wl_26 vdd gnd cell_6t
Xbit_r27_c49 bl_49 br_49 wl_27 vdd gnd cell_6t
Xbit_r28_c49 bl_49 br_49 wl_28 vdd gnd cell_6t
Xbit_r29_c49 bl_49 br_49 wl_29 vdd gnd cell_6t
Xbit_r30_c49 bl_49 br_49 wl_30 vdd gnd cell_6t
Xbit_r31_c49 bl_49 br_49 wl_31 vdd gnd cell_6t
Xbit_r32_c49 bl_49 br_49 wl_32 vdd gnd cell_6t
Xbit_r33_c49 bl_49 br_49 wl_33 vdd gnd cell_6t
Xbit_r34_c49 bl_49 br_49 wl_34 vdd gnd cell_6t
Xbit_r35_c49 bl_49 br_49 wl_35 vdd gnd cell_6t
Xbit_r36_c49 bl_49 br_49 wl_36 vdd gnd cell_6t
Xbit_r37_c49 bl_49 br_49 wl_37 vdd gnd cell_6t
Xbit_r38_c49 bl_49 br_49 wl_38 vdd gnd cell_6t
Xbit_r39_c49 bl_49 br_49 wl_39 vdd gnd cell_6t
Xbit_r40_c49 bl_49 br_49 wl_40 vdd gnd cell_6t
Xbit_r41_c49 bl_49 br_49 wl_41 vdd gnd cell_6t
Xbit_r42_c49 bl_49 br_49 wl_42 vdd gnd cell_6t
Xbit_r43_c49 bl_49 br_49 wl_43 vdd gnd cell_6t
Xbit_r44_c49 bl_49 br_49 wl_44 vdd gnd cell_6t
Xbit_r45_c49 bl_49 br_49 wl_45 vdd gnd cell_6t
Xbit_r46_c49 bl_49 br_49 wl_46 vdd gnd cell_6t
Xbit_r47_c49 bl_49 br_49 wl_47 vdd gnd cell_6t
Xbit_r48_c49 bl_49 br_49 wl_48 vdd gnd cell_6t
Xbit_r49_c49 bl_49 br_49 wl_49 vdd gnd cell_6t
Xbit_r50_c49 bl_49 br_49 wl_50 vdd gnd cell_6t
Xbit_r51_c49 bl_49 br_49 wl_51 vdd gnd cell_6t
Xbit_r52_c49 bl_49 br_49 wl_52 vdd gnd cell_6t
Xbit_r53_c49 bl_49 br_49 wl_53 vdd gnd cell_6t
Xbit_r54_c49 bl_49 br_49 wl_54 vdd gnd cell_6t
Xbit_r55_c49 bl_49 br_49 wl_55 vdd gnd cell_6t
Xbit_r56_c49 bl_49 br_49 wl_56 vdd gnd cell_6t
Xbit_r57_c49 bl_49 br_49 wl_57 vdd gnd cell_6t
Xbit_r58_c49 bl_49 br_49 wl_58 vdd gnd cell_6t
Xbit_r59_c49 bl_49 br_49 wl_59 vdd gnd cell_6t
Xbit_r60_c49 bl_49 br_49 wl_60 vdd gnd cell_6t
Xbit_r61_c49 bl_49 br_49 wl_61 vdd gnd cell_6t
Xbit_r62_c49 bl_49 br_49 wl_62 vdd gnd cell_6t
Xbit_r63_c49 bl_49 br_49 wl_63 vdd gnd cell_6t
Xbit_r64_c49 bl_49 br_49 wl_64 vdd gnd cell_6t
Xbit_r65_c49 bl_49 br_49 wl_65 vdd gnd cell_6t
Xbit_r66_c49 bl_49 br_49 wl_66 vdd gnd cell_6t
Xbit_r67_c49 bl_49 br_49 wl_67 vdd gnd cell_6t
Xbit_r68_c49 bl_49 br_49 wl_68 vdd gnd cell_6t
Xbit_r69_c49 bl_49 br_49 wl_69 vdd gnd cell_6t
Xbit_r70_c49 bl_49 br_49 wl_70 vdd gnd cell_6t
Xbit_r71_c49 bl_49 br_49 wl_71 vdd gnd cell_6t
Xbit_r72_c49 bl_49 br_49 wl_72 vdd gnd cell_6t
Xbit_r73_c49 bl_49 br_49 wl_73 vdd gnd cell_6t
Xbit_r74_c49 bl_49 br_49 wl_74 vdd gnd cell_6t
Xbit_r75_c49 bl_49 br_49 wl_75 vdd gnd cell_6t
Xbit_r76_c49 bl_49 br_49 wl_76 vdd gnd cell_6t
Xbit_r77_c49 bl_49 br_49 wl_77 vdd gnd cell_6t
Xbit_r78_c49 bl_49 br_49 wl_78 vdd gnd cell_6t
Xbit_r79_c49 bl_49 br_49 wl_79 vdd gnd cell_6t
Xbit_r80_c49 bl_49 br_49 wl_80 vdd gnd cell_6t
Xbit_r81_c49 bl_49 br_49 wl_81 vdd gnd cell_6t
Xbit_r82_c49 bl_49 br_49 wl_82 vdd gnd cell_6t
Xbit_r83_c49 bl_49 br_49 wl_83 vdd gnd cell_6t
Xbit_r84_c49 bl_49 br_49 wl_84 vdd gnd cell_6t
Xbit_r85_c49 bl_49 br_49 wl_85 vdd gnd cell_6t
Xbit_r86_c49 bl_49 br_49 wl_86 vdd gnd cell_6t
Xbit_r87_c49 bl_49 br_49 wl_87 vdd gnd cell_6t
Xbit_r88_c49 bl_49 br_49 wl_88 vdd gnd cell_6t
Xbit_r89_c49 bl_49 br_49 wl_89 vdd gnd cell_6t
Xbit_r90_c49 bl_49 br_49 wl_90 vdd gnd cell_6t
Xbit_r91_c49 bl_49 br_49 wl_91 vdd gnd cell_6t
Xbit_r92_c49 bl_49 br_49 wl_92 vdd gnd cell_6t
Xbit_r93_c49 bl_49 br_49 wl_93 vdd gnd cell_6t
Xbit_r94_c49 bl_49 br_49 wl_94 vdd gnd cell_6t
Xbit_r95_c49 bl_49 br_49 wl_95 vdd gnd cell_6t
Xbit_r96_c49 bl_49 br_49 wl_96 vdd gnd cell_6t
Xbit_r97_c49 bl_49 br_49 wl_97 vdd gnd cell_6t
Xbit_r98_c49 bl_49 br_49 wl_98 vdd gnd cell_6t
Xbit_r99_c49 bl_49 br_49 wl_99 vdd gnd cell_6t
Xbit_r100_c49 bl_49 br_49 wl_100 vdd gnd cell_6t
Xbit_r101_c49 bl_49 br_49 wl_101 vdd gnd cell_6t
Xbit_r102_c49 bl_49 br_49 wl_102 vdd gnd cell_6t
Xbit_r103_c49 bl_49 br_49 wl_103 vdd gnd cell_6t
Xbit_r104_c49 bl_49 br_49 wl_104 vdd gnd cell_6t
Xbit_r105_c49 bl_49 br_49 wl_105 vdd gnd cell_6t
Xbit_r106_c49 bl_49 br_49 wl_106 vdd gnd cell_6t
Xbit_r107_c49 bl_49 br_49 wl_107 vdd gnd cell_6t
Xbit_r108_c49 bl_49 br_49 wl_108 vdd gnd cell_6t
Xbit_r109_c49 bl_49 br_49 wl_109 vdd gnd cell_6t
Xbit_r110_c49 bl_49 br_49 wl_110 vdd gnd cell_6t
Xbit_r111_c49 bl_49 br_49 wl_111 vdd gnd cell_6t
Xbit_r112_c49 bl_49 br_49 wl_112 vdd gnd cell_6t
Xbit_r113_c49 bl_49 br_49 wl_113 vdd gnd cell_6t
Xbit_r114_c49 bl_49 br_49 wl_114 vdd gnd cell_6t
Xbit_r115_c49 bl_49 br_49 wl_115 vdd gnd cell_6t
Xbit_r116_c49 bl_49 br_49 wl_116 vdd gnd cell_6t
Xbit_r117_c49 bl_49 br_49 wl_117 vdd gnd cell_6t
Xbit_r118_c49 bl_49 br_49 wl_118 vdd gnd cell_6t
Xbit_r119_c49 bl_49 br_49 wl_119 vdd gnd cell_6t
Xbit_r120_c49 bl_49 br_49 wl_120 vdd gnd cell_6t
Xbit_r121_c49 bl_49 br_49 wl_121 vdd gnd cell_6t
Xbit_r122_c49 bl_49 br_49 wl_122 vdd gnd cell_6t
Xbit_r123_c49 bl_49 br_49 wl_123 vdd gnd cell_6t
Xbit_r124_c49 bl_49 br_49 wl_124 vdd gnd cell_6t
Xbit_r125_c49 bl_49 br_49 wl_125 vdd gnd cell_6t
Xbit_r126_c49 bl_49 br_49 wl_126 vdd gnd cell_6t
Xbit_r127_c49 bl_49 br_49 wl_127 vdd gnd cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd cell_6t
Xbit_r1_c50 bl_50 br_50 wl_1 vdd gnd cell_6t
Xbit_r2_c50 bl_50 br_50 wl_2 vdd gnd cell_6t
Xbit_r3_c50 bl_50 br_50 wl_3 vdd gnd cell_6t
Xbit_r4_c50 bl_50 br_50 wl_4 vdd gnd cell_6t
Xbit_r5_c50 bl_50 br_50 wl_5 vdd gnd cell_6t
Xbit_r6_c50 bl_50 br_50 wl_6 vdd gnd cell_6t
Xbit_r7_c50 bl_50 br_50 wl_7 vdd gnd cell_6t
Xbit_r8_c50 bl_50 br_50 wl_8 vdd gnd cell_6t
Xbit_r9_c50 bl_50 br_50 wl_9 vdd gnd cell_6t
Xbit_r10_c50 bl_50 br_50 wl_10 vdd gnd cell_6t
Xbit_r11_c50 bl_50 br_50 wl_11 vdd gnd cell_6t
Xbit_r12_c50 bl_50 br_50 wl_12 vdd gnd cell_6t
Xbit_r13_c50 bl_50 br_50 wl_13 vdd gnd cell_6t
Xbit_r14_c50 bl_50 br_50 wl_14 vdd gnd cell_6t
Xbit_r15_c50 bl_50 br_50 wl_15 vdd gnd cell_6t
Xbit_r16_c50 bl_50 br_50 wl_16 vdd gnd cell_6t
Xbit_r17_c50 bl_50 br_50 wl_17 vdd gnd cell_6t
Xbit_r18_c50 bl_50 br_50 wl_18 vdd gnd cell_6t
Xbit_r19_c50 bl_50 br_50 wl_19 vdd gnd cell_6t
Xbit_r20_c50 bl_50 br_50 wl_20 vdd gnd cell_6t
Xbit_r21_c50 bl_50 br_50 wl_21 vdd gnd cell_6t
Xbit_r22_c50 bl_50 br_50 wl_22 vdd gnd cell_6t
Xbit_r23_c50 bl_50 br_50 wl_23 vdd gnd cell_6t
Xbit_r24_c50 bl_50 br_50 wl_24 vdd gnd cell_6t
Xbit_r25_c50 bl_50 br_50 wl_25 vdd gnd cell_6t
Xbit_r26_c50 bl_50 br_50 wl_26 vdd gnd cell_6t
Xbit_r27_c50 bl_50 br_50 wl_27 vdd gnd cell_6t
Xbit_r28_c50 bl_50 br_50 wl_28 vdd gnd cell_6t
Xbit_r29_c50 bl_50 br_50 wl_29 vdd gnd cell_6t
Xbit_r30_c50 bl_50 br_50 wl_30 vdd gnd cell_6t
Xbit_r31_c50 bl_50 br_50 wl_31 vdd gnd cell_6t
Xbit_r32_c50 bl_50 br_50 wl_32 vdd gnd cell_6t
Xbit_r33_c50 bl_50 br_50 wl_33 vdd gnd cell_6t
Xbit_r34_c50 bl_50 br_50 wl_34 vdd gnd cell_6t
Xbit_r35_c50 bl_50 br_50 wl_35 vdd gnd cell_6t
Xbit_r36_c50 bl_50 br_50 wl_36 vdd gnd cell_6t
Xbit_r37_c50 bl_50 br_50 wl_37 vdd gnd cell_6t
Xbit_r38_c50 bl_50 br_50 wl_38 vdd gnd cell_6t
Xbit_r39_c50 bl_50 br_50 wl_39 vdd gnd cell_6t
Xbit_r40_c50 bl_50 br_50 wl_40 vdd gnd cell_6t
Xbit_r41_c50 bl_50 br_50 wl_41 vdd gnd cell_6t
Xbit_r42_c50 bl_50 br_50 wl_42 vdd gnd cell_6t
Xbit_r43_c50 bl_50 br_50 wl_43 vdd gnd cell_6t
Xbit_r44_c50 bl_50 br_50 wl_44 vdd gnd cell_6t
Xbit_r45_c50 bl_50 br_50 wl_45 vdd gnd cell_6t
Xbit_r46_c50 bl_50 br_50 wl_46 vdd gnd cell_6t
Xbit_r47_c50 bl_50 br_50 wl_47 vdd gnd cell_6t
Xbit_r48_c50 bl_50 br_50 wl_48 vdd gnd cell_6t
Xbit_r49_c50 bl_50 br_50 wl_49 vdd gnd cell_6t
Xbit_r50_c50 bl_50 br_50 wl_50 vdd gnd cell_6t
Xbit_r51_c50 bl_50 br_50 wl_51 vdd gnd cell_6t
Xbit_r52_c50 bl_50 br_50 wl_52 vdd gnd cell_6t
Xbit_r53_c50 bl_50 br_50 wl_53 vdd gnd cell_6t
Xbit_r54_c50 bl_50 br_50 wl_54 vdd gnd cell_6t
Xbit_r55_c50 bl_50 br_50 wl_55 vdd gnd cell_6t
Xbit_r56_c50 bl_50 br_50 wl_56 vdd gnd cell_6t
Xbit_r57_c50 bl_50 br_50 wl_57 vdd gnd cell_6t
Xbit_r58_c50 bl_50 br_50 wl_58 vdd gnd cell_6t
Xbit_r59_c50 bl_50 br_50 wl_59 vdd gnd cell_6t
Xbit_r60_c50 bl_50 br_50 wl_60 vdd gnd cell_6t
Xbit_r61_c50 bl_50 br_50 wl_61 vdd gnd cell_6t
Xbit_r62_c50 bl_50 br_50 wl_62 vdd gnd cell_6t
Xbit_r63_c50 bl_50 br_50 wl_63 vdd gnd cell_6t
Xbit_r64_c50 bl_50 br_50 wl_64 vdd gnd cell_6t
Xbit_r65_c50 bl_50 br_50 wl_65 vdd gnd cell_6t
Xbit_r66_c50 bl_50 br_50 wl_66 vdd gnd cell_6t
Xbit_r67_c50 bl_50 br_50 wl_67 vdd gnd cell_6t
Xbit_r68_c50 bl_50 br_50 wl_68 vdd gnd cell_6t
Xbit_r69_c50 bl_50 br_50 wl_69 vdd gnd cell_6t
Xbit_r70_c50 bl_50 br_50 wl_70 vdd gnd cell_6t
Xbit_r71_c50 bl_50 br_50 wl_71 vdd gnd cell_6t
Xbit_r72_c50 bl_50 br_50 wl_72 vdd gnd cell_6t
Xbit_r73_c50 bl_50 br_50 wl_73 vdd gnd cell_6t
Xbit_r74_c50 bl_50 br_50 wl_74 vdd gnd cell_6t
Xbit_r75_c50 bl_50 br_50 wl_75 vdd gnd cell_6t
Xbit_r76_c50 bl_50 br_50 wl_76 vdd gnd cell_6t
Xbit_r77_c50 bl_50 br_50 wl_77 vdd gnd cell_6t
Xbit_r78_c50 bl_50 br_50 wl_78 vdd gnd cell_6t
Xbit_r79_c50 bl_50 br_50 wl_79 vdd gnd cell_6t
Xbit_r80_c50 bl_50 br_50 wl_80 vdd gnd cell_6t
Xbit_r81_c50 bl_50 br_50 wl_81 vdd gnd cell_6t
Xbit_r82_c50 bl_50 br_50 wl_82 vdd gnd cell_6t
Xbit_r83_c50 bl_50 br_50 wl_83 vdd gnd cell_6t
Xbit_r84_c50 bl_50 br_50 wl_84 vdd gnd cell_6t
Xbit_r85_c50 bl_50 br_50 wl_85 vdd gnd cell_6t
Xbit_r86_c50 bl_50 br_50 wl_86 vdd gnd cell_6t
Xbit_r87_c50 bl_50 br_50 wl_87 vdd gnd cell_6t
Xbit_r88_c50 bl_50 br_50 wl_88 vdd gnd cell_6t
Xbit_r89_c50 bl_50 br_50 wl_89 vdd gnd cell_6t
Xbit_r90_c50 bl_50 br_50 wl_90 vdd gnd cell_6t
Xbit_r91_c50 bl_50 br_50 wl_91 vdd gnd cell_6t
Xbit_r92_c50 bl_50 br_50 wl_92 vdd gnd cell_6t
Xbit_r93_c50 bl_50 br_50 wl_93 vdd gnd cell_6t
Xbit_r94_c50 bl_50 br_50 wl_94 vdd gnd cell_6t
Xbit_r95_c50 bl_50 br_50 wl_95 vdd gnd cell_6t
Xbit_r96_c50 bl_50 br_50 wl_96 vdd gnd cell_6t
Xbit_r97_c50 bl_50 br_50 wl_97 vdd gnd cell_6t
Xbit_r98_c50 bl_50 br_50 wl_98 vdd gnd cell_6t
Xbit_r99_c50 bl_50 br_50 wl_99 vdd gnd cell_6t
Xbit_r100_c50 bl_50 br_50 wl_100 vdd gnd cell_6t
Xbit_r101_c50 bl_50 br_50 wl_101 vdd gnd cell_6t
Xbit_r102_c50 bl_50 br_50 wl_102 vdd gnd cell_6t
Xbit_r103_c50 bl_50 br_50 wl_103 vdd gnd cell_6t
Xbit_r104_c50 bl_50 br_50 wl_104 vdd gnd cell_6t
Xbit_r105_c50 bl_50 br_50 wl_105 vdd gnd cell_6t
Xbit_r106_c50 bl_50 br_50 wl_106 vdd gnd cell_6t
Xbit_r107_c50 bl_50 br_50 wl_107 vdd gnd cell_6t
Xbit_r108_c50 bl_50 br_50 wl_108 vdd gnd cell_6t
Xbit_r109_c50 bl_50 br_50 wl_109 vdd gnd cell_6t
Xbit_r110_c50 bl_50 br_50 wl_110 vdd gnd cell_6t
Xbit_r111_c50 bl_50 br_50 wl_111 vdd gnd cell_6t
Xbit_r112_c50 bl_50 br_50 wl_112 vdd gnd cell_6t
Xbit_r113_c50 bl_50 br_50 wl_113 vdd gnd cell_6t
Xbit_r114_c50 bl_50 br_50 wl_114 vdd gnd cell_6t
Xbit_r115_c50 bl_50 br_50 wl_115 vdd gnd cell_6t
Xbit_r116_c50 bl_50 br_50 wl_116 vdd gnd cell_6t
Xbit_r117_c50 bl_50 br_50 wl_117 vdd gnd cell_6t
Xbit_r118_c50 bl_50 br_50 wl_118 vdd gnd cell_6t
Xbit_r119_c50 bl_50 br_50 wl_119 vdd gnd cell_6t
Xbit_r120_c50 bl_50 br_50 wl_120 vdd gnd cell_6t
Xbit_r121_c50 bl_50 br_50 wl_121 vdd gnd cell_6t
Xbit_r122_c50 bl_50 br_50 wl_122 vdd gnd cell_6t
Xbit_r123_c50 bl_50 br_50 wl_123 vdd gnd cell_6t
Xbit_r124_c50 bl_50 br_50 wl_124 vdd gnd cell_6t
Xbit_r125_c50 bl_50 br_50 wl_125 vdd gnd cell_6t
Xbit_r126_c50 bl_50 br_50 wl_126 vdd gnd cell_6t
Xbit_r127_c50 bl_50 br_50 wl_127 vdd gnd cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd cell_6t
Xbit_r1_c51 bl_51 br_51 wl_1 vdd gnd cell_6t
Xbit_r2_c51 bl_51 br_51 wl_2 vdd gnd cell_6t
Xbit_r3_c51 bl_51 br_51 wl_3 vdd gnd cell_6t
Xbit_r4_c51 bl_51 br_51 wl_4 vdd gnd cell_6t
Xbit_r5_c51 bl_51 br_51 wl_5 vdd gnd cell_6t
Xbit_r6_c51 bl_51 br_51 wl_6 vdd gnd cell_6t
Xbit_r7_c51 bl_51 br_51 wl_7 vdd gnd cell_6t
Xbit_r8_c51 bl_51 br_51 wl_8 vdd gnd cell_6t
Xbit_r9_c51 bl_51 br_51 wl_9 vdd gnd cell_6t
Xbit_r10_c51 bl_51 br_51 wl_10 vdd gnd cell_6t
Xbit_r11_c51 bl_51 br_51 wl_11 vdd gnd cell_6t
Xbit_r12_c51 bl_51 br_51 wl_12 vdd gnd cell_6t
Xbit_r13_c51 bl_51 br_51 wl_13 vdd gnd cell_6t
Xbit_r14_c51 bl_51 br_51 wl_14 vdd gnd cell_6t
Xbit_r15_c51 bl_51 br_51 wl_15 vdd gnd cell_6t
Xbit_r16_c51 bl_51 br_51 wl_16 vdd gnd cell_6t
Xbit_r17_c51 bl_51 br_51 wl_17 vdd gnd cell_6t
Xbit_r18_c51 bl_51 br_51 wl_18 vdd gnd cell_6t
Xbit_r19_c51 bl_51 br_51 wl_19 vdd gnd cell_6t
Xbit_r20_c51 bl_51 br_51 wl_20 vdd gnd cell_6t
Xbit_r21_c51 bl_51 br_51 wl_21 vdd gnd cell_6t
Xbit_r22_c51 bl_51 br_51 wl_22 vdd gnd cell_6t
Xbit_r23_c51 bl_51 br_51 wl_23 vdd gnd cell_6t
Xbit_r24_c51 bl_51 br_51 wl_24 vdd gnd cell_6t
Xbit_r25_c51 bl_51 br_51 wl_25 vdd gnd cell_6t
Xbit_r26_c51 bl_51 br_51 wl_26 vdd gnd cell_6t
Xbit_r27_c51 bl_51 br_51 wl_27 vdd gnd cell_6t
Xbit_r28_c51 bl_51 br_51 wl_28 vdd gnd cell_6t
Xbit_r29_c51 bl_51 br_51 wl_29 vdd gnd cell_6t
Xbit_r30_c51 bl_51 br_51 wl_30 vdd gnd cell_6t
Xbit_r31_c51 bl_51 br_51 wl_31 vdd gnd cell_6t
Xbit_r32_c51 bl_51 br_51 wl_32 vdd gnd cell_6t
Xbit_r33_c51 bl_51 br_51 wl_33 vdd gnd cell_6t
Xbit_r34_c51 bl_51 br_51 wl_34 vdd gnd cell_6t
Xbit_r35_c51 bl_51 br_51 wl_35 vdd gnd cell_6t
Xbit_r36_c51 bl_51 br_51 wl_36 vdd gnd cell_6t
Xbit_r37_c51 bl_51 br_51 wl_37 vdd gnd cell_6t
Xbit_r38_c51 bl_51 br_51 wl_38 vdd gnd cell_6t
Xbit_r39_c51 bl_51 br_51 wl_39 vdd gnd cell_6t
Xbit_r40_c51 bl_51 br_51 wl_40 vdd gnd cell_6t
Xbit_r41_c51 bl_51 br_51 wl_41 vdd gnd cell_6t
Xbit_r42_c51 bl_51 br_51 wl_42 vdd gnd cell_6t
Xbit_r43_c51 bl_51 br_51 wl_43 vdd gnd cell_6t
Xbit_r44_c51 bl_51 br_51 wl_44 vdd gnd cell_6t
Xbit_r45_c51 bl_51 br_51 wl_45 vdd gnd cell_6t
Xbit_r46_c51 bl_51 br_51 wl_46 vdd gnd cell_6t
Xbit_r47_c51 bl_51 br_51 wl_47 vdd gnd cell_6t
Xbit_r48_c51 bl_51 br_51 wl_48 vdd gnd cell_6t
Xbit_r49_c51 bl_51 br_51 wl_49 vdd gnd cell_6t
Xbit_r50_c51 bl_51 br_51 wl_50 vdd gnd cell_6t
Xbit_r51_c51 bl_51 br_51 wl_51 vdd gnd cell_6t
Xbit_r52_c51 bl_51 br_51 wl_52 vdd gnd cell_6t
Xbit_r53_c51 bl_51 br_51 wl_53 vdd gnd cell_6t
Xbit_r54_c51 bl_51 br_51 wl_54 vdd gnd cell_6t
Xbit_r55_c51 bl_51 br_51 wl_55 vdd gnd cell_6t
Xbit_r56_c51 bl_51 br_51 wl_56 vdd gnd cell_6t
Xbit_r57_c51 bl_51 br_51 wl_57 vdd gnd cell_6t
Xbit_r58_c51 bl_51 br_51 wl_58 vdd gnd cell_6t
Xbit_r59_c51 bl_51 br_51 wl_59 vdd gnd cell_6t
Xbit_r60_c51 bl_51 br_51 wl_60 vdd gnd cell_6t
Xbit_r61_c51 bl_51 br_51 wl_61 vdd gnd cell_6t
Xbit_r62_c51 bl_51 br_51 wl_62 vdd gnd cell_6t
Xbit_r63_c51 bl_51 br_51 wl_63 vdd gnd cell_6t
Xbit_r64_c51 bl_51 br_51 wl_64 vdd gnd cell_6t
Xbit_r65_c51 bl_51 br_51 wl_65 vdd gnd cell_6t
Xbit_r66_c51 bl_51 br_51 wl_66 vdd gnd cell_6t
Xbit_r67_c51 bl_51 br_51 wl_67 vdd gnd cell_6t
Xbit_r68_c51 bl_51 br_51 wl_68 vdd gnd cell_6t
Xbit_r69_c51 bl_51 br_51 wl_69 vdd gnd cell_6t
Xbit_r70_c51 bl_51 br_51 wl_70 vdd gnd cell_6t
Xbit_r71_c51 bl_51 br_51 wl_71 vdd gnd cell_6t
Xbit_r72_c51 bl_51 br_51 wl_72 vdd gnd cell_6t
Xbit_r73_c51 bl_51 br_51 wl_73 vdd gnd cell_6t
Xbit_r74_c51 bl_51 br_51 wl_74 vdd gnd cell_6t
Xbit_r75_c51 bl_51 br_51 wl_75 vdd gnd cell_6t
Xbit_r76_c51 bl_51 br_51 wl_76 vdd gnd cell_6t
Xbit_r77_c51 bl_51 br_51 wl_77 vdd gnd cell_6t
Xbit_r78_c51 bl_51 br_51 wl_78 vdd gnd cell_6t
Xbit_r79_c51 bl_51 br_51 wl_79 vdd gnd cell_6t
Xbit_r80_c51 bl_51 br_51 wl_80 vdd gnd cell_6t
Xbit_r81_c51 bl_51 br_51 wl_81 vdd gnd cell_6t
Xbit_r82_c51 bl_51 br_51 wl_82 vdd gnd cell_6t
Xbit_r83_c51 bl_51 br_51 wl_83 vdd gnd cell_6t
Xbit_r84_c51 bl_51 br_51 wl_84 vdd gnd cell_6t
Xbit_r85_c51 bl_51 br_51 wl_85 vdd gnd cell_6t
Xbit_r86_c51 bl_51 br_51 wl_86 vdd gnd cell_6t
Xbit_r87_c51 bl_51 br_51 wl_87 vdd gnd cell_6t
Xbit_r88_c51 bl_51 br_51 wl_88 vdd gnd cell_6t
Xbit_r89_c51 bl_51 br_51 wl_89 vdd gnd cell_6t
Xbit_r90_c51 bl_51 br_51 wl_90 vdd gnd cell_6t
Xbit_r91_c51 bl_51 br_51 wl_91 vdd gnd cell_6t
Xbit_r92_c51 bl_51 br_51 wl_92 vdd gnd cell_6t
Xbit_r93_c51 bl_51 br_51 wl_93 vdd gnd cell_6t
Xbit_r94_c51 bl_51 br_51 wl_94 vdd gnd cell_6t
Xbit_r95_c51 bl_51 br_51 wl_95 vdd gnd cell_6t
Xbit_r96_c51 bl_51 br_51 wl_96 vdd gnd cell_6t
Xbit_r97_c51 bl_51 br_51 wl_97 vdd gnd cell_6t
Xbit_r98_c51 bl_51 br_51 wl_98 vdd gnd cell_6t
Xbit_r99_c51 bl_51 br_51 wl_99 vdd gnd cell_6t
Xbit_r100_c51 bl_51 br_51 wl_100 vdd gnd cell_6t
Xbit_r101_c51 bl_51 br_51 wl_101 vdd gnd cell_6t
Xbit_r102_c51 bl_51 br_51 wl_102 vdd gnd cell_6t
Xbit_r103_c51 bl_51 br_51 wl_103 vdd gnd cell_6t
Xbit_r104_c51 bl_51 br_51 wl_104 vdd gnd cell_6t
Xbit_r105_c51 bl_51 br_51 wl_105 vdd gnd cell_6t
Xbit_r106_c51 bl_51 br_51 wl_106 vdd gnd cell_6t
Xbit_r107_c51 bl_51 br_51 wl_107 vdd gnd cell_6t
Xbit_r108_c51 bl_51 br_51 wl_108 vdd gnd cell_6t
Xbit_r109_c51 bl_51 br_51 wl_109 vdd gnd cell_6t
Xbit_r110_c51 bl_51 br_51 wl_110 vdd gnd cell_6t
Xbit_r111_c51 bl_51 br_51 wl_111 vdd gnd cell_6t
Xbit_r112_c51 bl_51 br_51 wl_112 vdd gnd cell_6t
Xbit_r113_c51 bl_51 br_51 wl_113 vdd gnd cell_6t
Xbit_r114_c51 bl_51 br_51 wl_114 vdd gnd cell_6t
Xbit_r115_c51 bl_51 br_51 wl_115 vdd gnd cell_6t
Xbit_r116_c51 bl_51 br_51 wl_116 vdd gnd cell_6t
Xbit_r117_c51 bl_51 br_51 wl_117 vdd gnd cell_6t
Xbit_r118_c51 bl_51 br_51 wl_118 vdd gnd cell_6t
Xbit_r119_c51 bl_51 br_51 wl_119 vdd gnd cell_6t
Xbit_r120_c51 bl_51 br_51 wl_120 vdd gnd cell_6t
Xbit_r121_c51 bl_51 br_51 wl_121 vdd gnd cell_6t
Xbit_r122_c51 bl_51 br_51 wl_122 vdd gnd cell_6t
Xbit_r123_c51 bl_51 br_51 wl_123 vdd gnd cell_6t
Xbit_r124_c51 bl_51 br_51 wl_124 vdd gnd cell_6t
Xbit_r125_c51 bl_51 br_51 wl_125 vdd gnd cell_6t
Xbit_r126_c51 bl_51 br_51 wl_126 vdd gnd cell_6t
Xbit_r127_c51 bl_51 br_51 wl_127 vdd gnd cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd cell_6t
Xbit_r1_c52 bl_52 br_52 wl_1 vdd gnd cell_6t
Xbit_r2_c52 bl_52 br_52 wl_2 vdd gnd cell_6t
Xbit_r3_c52 bl_52 br_52 wl_3 vdd gnd cell_6t
Xbit_r4_c52 bl_52 br_52 wl_4 vdd gnd cell_6t
Xbit_r5_c52 bl_52 br_52 wl_5 vdd gnd cell_6t
Xbit_r6_c52 bl_52 br_52 wl_6 vdd gnd cell_6t
Xbit_r7_c52 bl_52 br_52 wl_7 vdd gnd cell_6t
Xbit_r8_c52 bl_52 br_52 wl_8 vdd gnd cell_6t
Xbit_r9_c52 bl_52 br_52 wl_9 vdd gnd cell_6t
Xbit_r10_c52 bl_52 br_52 wl_10 vdd gnd cell_6t
Xbit_r11_c52 bl_52 br_52 wl_11 vdd gnd cell_6t
Xbit_r12_c52 bl_52 br_52 wl_12 vdd gnd cell_6t
Xbit_r13_c52 bl_52 br_52 wl_13 vdd gnd cell_6t
Xbit_r14_c52 bl_52 br_52 wl_14 vdd gnd cell_6t
Xbit_r15_c52 bl_52 br_52 wl_15 vdd gnd cell_6t
Xbit_r16_c52 bl_52 br_52 wl_16 vdd gnd cell_6t
Xbit_r17_c52 bl_52 br_52 wl_17 vdd gnd cell_6t
Xbit_r18_c52 bl_52 br_52 wl_18 vdd gnd cell_6t
Xbit_r19_c52 bl_52 br_52 wl_19 vdd gnd cell_6t
Xbit_r20_c52 bl_52 br_52 wl_20 vdd gnd cell_6t
Xbit_r21_c52 bl_52 br_52 wl_21 vdd gnd cell_6t
Xbit_r22_c52 bl_52 br_52 wl_22 vdd gnd cell_6t
Xbit_r23_c52 bl_52 br_52 wl_23 vdd gnd cell_6t
Xbit_r24_c52 bl_52 br_52 wl_24 vdd gnd cell_6t
Xbit_r25_c52 bl_52 br_52 wl_25 vdd gnd cell_6t
Xbit_r26_c52 bl_52 br_52 wl_26 vdd gnd cell_6t
Xbit_r27_c52 bl_52 br_52 wl_27 vdd gnd cell_6t
Xbit_r28_c52 bl_52 br_52 wl_28 vdd gnd cell_6t
Xbit_r29_c52 bl_52 br_52 wl_29 vdd gnd cell_6t
Xbit_r30_c52 bl_52 br_52 wl_30 vdd gnd cell_6t
Xbit_r31_c52 bl_52 br_52 wl_31 vdd gnd cell_6t
Xbit_r32_c52 bl_52 br_52 wl_32 vdd gnd cell_6t
Xbit_r33_c52 bl_52 br_52 wl_33 vdd gnd cell_6t
Xbit_r34_c52 bl_52 br_52 wl_34 vdd gnd cell_6t
Xbit_r35_c52 bl_52 br_52 wl_35 vdd gnd cell_6t
Xbit_r36_c52 bl_52 br_52 wl_36 vdd gnd cell_6t
Xbit_r37_c52 bl_52 br_52 wl_37 vdd gnd cell_6t
Xbit_r38_c52 bl_52 br_52 wl_38 vdd gnd cell_6t
Xbit_r39_c52 bl_52 br_52 wl_39 vdd gnd cell_6t
Xbit_r40_c52 bl_52 br_52 wl_40 vdd gnd cell_6t
Xbit_r41_c52 bl_52 br_52 wl_41 vdd gnd cell_6t
Xbit_r42_c52 bl_52 br_52 wl_42 vdd gnd cell_6t
Xbit_r43_c52 bl_52 br_52 wl_43 vdd gnd cell_6t
Xbit_r44_c52 bl_52 br_52 wl_44 vdd gnd cell_6t
Xbit_r45_c52 bl_52 br_52 wl_45 vdd gnd cell_6t
Xbit_r46_c52 bl_52 br_52 wl_46 vdd gnd cell_6t
Xbit_r47_c52 bl_52 br_52 wl_47 vdd gnd cell_6t
Xbit_r48_c52 bl_52 br_52 wl_48 vdd gnd cell_6t
Xbit_r49_c52 bl_52 br_52 wl_49 vdd gnd cell_6t
Xbit_r50_c52 bl_52 br_52 wl_50 vdd gnd cell_6t
Xbit_r51_c52 bl_52 br_52 wl_51 vdd gnd cell_6t
Xbit_r52_c52 bl_52 br_52 wl_52 vdd gnd cell_6t
Xbit_r53_c52 bl_52 br_52 wl_53 vdd gnd cell_6t
Xbit_r54_c52 bl_52 br_52 wl_54 vdd gnd cell_6t
Xbit_r55_c52 bl_52 br_52 wl_55 vdd gnd cell_6t
Xbit_r56_c52 bl_52 br_52 wl_56 vdd gnd cell_6t
Xbit_r57_c52 bl_52 br_52 wl_57 vdd gnd cell_6t
Xbit_r58_c52 bl_52 br_52 wl_58 vdd gnd cell_6t
Xbit_r59_c52 bl_52 br_52 wl_59 vdd gnd cell_6t
Xbit_r60_c52 bl_52 br_52 wl_60 vdd gnd cell_6t
Xbit_r61_c52 bl_52 br_52 wl_61 vdd gnd cell_6t
Xbit_r62_c52 bl_52 br_52 wl_62 vdd gnd cell_6t
Xbit_r63_c52 bl_52 br_52 wl_63 vdd gnd cell_6t
Xbit_r64_c52 bl_52 br_52 wl_64 vdd gnd cell_6t
Xbit_r65_c52 bl_52 br_52 wl_65 vdd gnd cell_6t
Xbit_r66_c52 bl_52 br_52 wl_66 vdd gnd cell_6t
Xbit_r67_c52 bl_52 br_52 wl_67 vdd gnd cell_6t
Xbit_r68_c52 bl_52 br_52 wl_68 vdd gnd cell_6t
Xbit_r69_c52 bl_52 br_52 wl_69 vdd gnd cell_6t
Xbit_r70_c52 bl_52 br_52 wl_70 vdd gnd cell_6t
Xbit_r71_c52 bl_52 br_52 wl_71 vdd gnd cell_6t
Xbit_r72_c52 bl_52 br_52 wl_72 vdd gnd cell_6t
Xbit_r73_c52 bl_52 br_52 wl_73 vdd gnd cell_6t
Xbit_r74_c52 bl_52 br_52 wl_74 vdd gnd cell_6t
Xbit_r75_c52 bl_52 br_52 wl_75 vdd gnd cell_6t
Xbit_r76_c52 bl_52 br_52 wl_76 vdd gnd cell_6t
Xbit_r77_c52 bl_52 br_52 wl_77 vdd gnd cell_6t
Xbit_r78_c52 bl_52 br_52 wl_78 vdd gnd cell_6t
Xbit_r79_c52 bl_52 br_52 wl_79 vdd gnd cell_6t
Xbit_r80_c52 bl_52 br_52 wl_80 vdd gnd cell_6t
Xbit_r81_c52 bl_52 br_52 wl_81 vdd gnd cell_6t
Xbit_r82_c52 bl_52 br_52 wl_82 vdd gnd cell_6t
Xbit_r83_c52 bl_52 br_52 wl_83 vdd gnd cell_6t
Xbit_r84_c52 bl_52 br_52 wl_84 vdd gnd cell_6t
Xbit_r85_c52 bl_52 br_52 wl_85 vdd gnd cell_6t
Xbit_r86_c52 bl_52 br_52 wl_86 vdd gnd cell_6t
Xbit_r87_c52 bl_52 br_52 wl_87 vdd gnd cell_6t
Xbit_r88_c52 bl_52 br_52 wl_88 vdd gnd cell_6t
Xbit_r89_c52 bl_52 br_52 wl_89 vdd gnd cell_6t
Xbit_r90_c52 bl_52 br_52 wl_90 vdd gnd cell_6t
Xbit_r91_c52 bl_52 br_52 wl_91 vdd gnd cell_6t
Xbit_r92_c52 bl_52 br_52 wl_92 vdd gnd cell_6t
Xbit_r93_c52 bl_52 br_52 wl_93 vdd gnd cell_6t
Xbit_r94_c52 bl_52 br_52 wl_94 vdd gnd cell_6t
Xbit_r95_c52 bl_52 br_52 wl_95 vdd gnd cell_6t
Xbit_r96_c52 bl_52 br_52 wl_96 vdd gnd cell_6t
Xbit_r97_c52 bl_52 br_52 wl_97 vdd gnd cell_6t
Xbit_r98_c52 bl_52 br_52 wl_98 vdd gnd cell_6t
Xbit_r99_c52 bl_52 br_52 wl_99 vdd gnd cell_6t
Xbit_r100_c52 bl_52 br_52 wl_100 vdd gnd cell_6t
Xbit_r101_c52 bl_52 br_52 wl_101 vdd gnd cell_6t
Xbit_r102_c52 bl_52 br_52 wl_102 vdd gnd cell_6t
Xbit_r103_c52 bl_52 br_52 wl_103 vdd gnd cell_6t
Xbit_r104_c52 bl_52 br_52 wl_104 vdd gnd cell_6t
Xbit_r105_c52 bl_52 br_52 wl_105 vdd gnd cell_6t
Xbit_r106_c52 bl_52 br_52 wl_106 vdd gnd cell_6t
Xbit_r107_c52 bl_52 br_52 wl_107 vdd gnd cell_6t
Xbit_r108_c52 bl_52 br_52 wl_108 vdd gnd cell_6t
Xbit_r109_c52 bl_52 br_52 wl_109 vdd gnd cell_6t
Xbit_r110_c52 bl_52 br_52 wl_110 vdd gnd cell_6t
Xbit_r111_c52 bl_52 br_52 wl_111 vdd gnd cell_6t
Xbit_r112_c52 bl_52 br_52 wl_112 vdd gnd cell_6t
Xbit_r113_c52 bl_52 br_52 wl_113 vdd gnd cell_6t
Xbit_r114_c52 bl_52 br_52 wl_114 vdd gnd cell_6t
Xbit_r115_c52 bl_52 br_52 wl_115 vdd gnd cell_6t
Xbit_r116_c52 bl_52 br_52 wl_116 vdd gnd cell_6t
Xbit_r117_c52 bl_52 br_52 wl_117 vdd gnd cell_6t
Xbit_r118_c52 bl_52 br_52 wl_118 vdd gnd cell_6t
Xbit_r119_c52 bl_52 br_52 wl_119 vdd gnd cell_6t
Xbit_r120_c52 bl_52 br_52 wl_120 vdd gnd cell_6t
Xbit_r121_c52 bl_52 br_52 wl_121 vdd gnd cell_6t
Xbit_r122_c52 bl_52 br_52 wl_122 vdd gnd cell_6t
Xbit_r123_c52 bl_52 br_52 wl_123 vdd gnd cell_6t
Xbit_r124_c52 bl_52 br_52 wl_124 vdd gnd cell_6t
Xbit_r125_c52 bl_52 br_52 wl_125 vdd gnd cell_6t
Xbit_r126_c52 bl_52 br_52 wl_126 vdd gnd cell_6t
Xbit_r127_c52 bl_52 br_52 wl_127 vdd gnd cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd cell_6t
Xbit_r1_c53 bl_53 br_53 wl_1 vdd gnd cell_6t
Xbit_r2_c53 bl_53 br_53 wl_2 vdd gnd cell_6t
Xbit_r3_c53 bl_53 br_53 wl_3 vdd gnd cell_6t
Xbit_r4_c53 bl_53 br_53 wl_4 vdd gnd cell_6t
Xbit_r5_c53 bl_53 br_53 wl_5 vdd gnd cell_6t
Xbit_r6_c53 bl_53 br_53 wl_6 vdd gnd cell_6t
Xbit_r7_c53 bl_53 br_53 wl_7 vdd gnd cell_6t
Xbit_r8_c53 bl_53 br_53 wl_8 vdd gnd cell_6t
Xbit_r9_c53 bl_53 br_53 wl_9 vdd gnd cell_6t
Xbit_r10_c53 bl_53 br_53 wl_10 vdd gnd cell_6t
Xbit_r11_c53 bl_53 br_53 wl_11 vdd gnd cell_6t
Xbit_r12_c53 bl_53 br_53 wl_12 vdd gnd cell_6t
Xbit_r13_c53 bl_53 br_53 wl_13 vdd gnd cell_6t
Xbit_r14_c53 bl_53 br_53 wl_14 vdd gnd cell_6t
Xbit_r15_c53 bl_53 br_53 wl_15 vdd gnd cell_6t
Xbit_r16_c53 bl_53 br_53 wl_16 vdd gnd cell_6t
Xbit_r17_c53 bl_53 br_53 wl_17 vdd gnd cell_6t
Xbit_r18_c53 bl_53 br_53 wl_18 vdd gnd cell_6t
Xbit_r19_c53 bl_53 br_53 wl_19 vdd gnd cell_6t
Xbit_r20_c53 bl_53 br_53 wl_20 vdd gnd cell_6t
Xbit_r21_c53 bl_53 br_53 wl_21 vdd gnd cell_6t
Xbit_r22_c53 bl_53 br_53 wl_22 vdd gnd cell_6t
Xbit_r23_c53 bl_53 br_53 wl_23 vdd gnd cell_6t
Xbit_r24_c53 bl_53 br_53 wl_24 vdd gnd cell_6t
Xbit_r25_c53 bl_53 br_53 wl_25 vdd gnd cell_6t
Xbit_r26_c53 bl_53 br_53 wl_26 vdd gnd cell_6t
Xbit_r27_c53 bl_53 br_53 wl_27 vdd gnd cell_6t
Xbit_r28_c53 bl_53 br_53 wl_28 vdd gnd cell_6t
Xbit_r29_c53 bl_53 br_53 wl_29 vdd gnd cell_6t
Xbit_r30_c53 bl_53 br_53 wl_30 vdd gnd cell_6t
Xbit_r31_c53 bl_53 br_53 wl_31 vdd gnd cell_6t
Xbit_r32_c53 bl_53 br_53 wl_32 vdd gnd cell_6t
Xbit_r33_c53 bl_53 br_53 wl_33 vdd gnd cell_6t
Xbit_r34_c53 bl_53 br_53 wl_34 vdd gnd cell_6t
Xbit_r35_c53 bl_53 br_53 wl_35 vdd gnd cell_6t
Xbit_r36_c53 bl_53 br_53 wl_36 vdd gnd cell_6t
Xbit_r37_c53 bl_53 br_53 wl_37 vdd gnd cell_6t
Xbit_r38_c53 bl_53 br_53 wl_38 vdd gnd cell_6t
Xbit_r39_c53 bl_53 br_53 wl_39 vdd gnd cell_6t
Xbit_r40_c53 bl_53 br_53 wl_40 vdd gnd cell_6t
Xbit_r41_c53 bl_53 br_53 wl_41 vdd gnd cell_6t
Xbit_r42_c53 bl_53 br_53 wl_42 vdd gnd cell_6t
Xbit_r43_c53 bl_53 br_53 wl_43 vdd gnd cell_6t
Xbit_r44_c53 bl_53 br_53 wl_44 vdd gnd cell_6t
Xbit_r45_c53 bl_53 br_53 wl_45 vdd gnd cell_6t
Xbit_r46_c53 bl_53 br_53 wl_46 vdd gnd cell_6t
Xbit_r47_c53 bl_53 br_53 wl_47 vdd gnd cell_6t
Xbit_r48_c53 bl_53 br_53 wl_48 vdd gnd cell_6t
Xbit_r49_c53 bl_53 br_53 wl_49 vdd gnd cell_6t
Xbit_r50_c53 bl_53 br_53 wl_50 vdd gnd cell_6t
Xbit_r51_c53 bl_53 br_53 wl_51 vdd gnd cell_6t
Xbit_r52_c53 bl_53 br_53 wl_52 vdd gnd cell_6t
Xbit_r53_c53 bl_53 br_53 wl_53 vdd gnd cell_6t
Xbit_r54_c53 bl_53 br_53 wl_54 vdd gnd cell_6t
Xbit_r55_c53 bl_53 br_53 wl_55 vdd gnd cell_6t
Xbit_r56_c53 bl_53 br_53 wl_56 vdd gnd cell_6t
Xbit_r57_c53 bl_53 br_53 wl_57 vdd gnd cell_6t
Xbit_r58_c53 bl_53 br_53 wl_58 vdd gnd cell_6t
Xbit_r59_c53 bl_53 br_53 wl_59 vdd gnd cell_6t
Xbit_r60_c53 bl_53 br_53 wl_60 vdd gnd cell_6t
Xbit_r61_c53 bl_53 br_53 wl_61 vdd gnd cell_6t
Xbit_r62_c53 bl_53 br_53 wl_62 vdd gnd cell_6t
Xbit_r63_c53 bl_53 br_53 wl_63 vdd gnd cell_6t
Xbit_r64_c53 bl_53 br_53 wl_64 vdd gnd cell_6t
Xbit_r65_c53 bl_53 br_53 wl_65 vdd gnd cell_6t
Xbit_r66_c53 bl_53 br_53 wl_66 vdd gnd cell_6t
Xbit_r67_c53 bl_53 br_53 wl_67 vdd gnd cell_6t
Xbit_r68_c53 bl_53 br_53 wl_68 vdd gnd cell_6t
Xbit_r69_c53 bl_53 br_53 wl_69 vdd gnd cell_6t
Xbit_r70_c53 bl_53 br_53 wl_70 vdd gnd cell_6t
Xbit_r71_c53 bl_53 br_53 wl_71 vdd gnd cell_6t
Xbit_r72_c53 bl_53 br_53 wl_72 vdd gnd cell_6t
Xbit_r73_c53 bl_53 br_53 wl_73 vdd gnd cell_6t
Xbit_r74_c53 bl_53 br_53 wl_74 vdd gnd cell_6t
Xbit_r75_c53 bl_53 br_53 wl_75 vdd gnd cell_6t
Xbit_r76_c53 bl_53 br_53 wl_76 vdd gnd cell_6t
Xbit_r77_c53 bl_53 br_53 wl_77 vdd gnd cell_6t
Xbit_r78_c53 bl_53 br_53 wl_78 vdd gnd cell_6t
Xbit_r79_c53 bl_53 br_53 wl_79 vdd gnd cell_6t
Xbit_r80_c53 bl_53 br_53 wl_80 vdd gnd cell_6t
Xbit_r81_c53 bl_53 br_53 wl_81 vdd gnd cell_6t
Xbit_r82_c53 bl_53 br_53 wl_82 vdd gnd cell_6t
Xbit_r83_c53 bl_53 br_53 wl_83 vdd gnd cell_6t
Xbit_r84_c53 bl_53 br_53 wl_84 vdd gnd cell_6t
Xbit_r85_c53 bl_53 br_53 wl_85 vdd gnd cell_6t
Xbit_r86_c53 bl_53 br_53 wl_86 vdd gnd cell_6t
Xbit_r87_c53 bl_53 br_53 wl_87 vdd gnd cell_6t
Xbit_r88_c53 bl_53 br_53 wl_88 vdd gnd cell_6t
Xbit_r89_c53 bl_53 br_53 wl_89 vdd gnd cell_6t
Xbit_r90_c53 bl_53 br_53 wl_90 vdd gnd cell_6t
Xbit_r91_c53 bl_53 br_53 wl_91 vdd gnd cell_6t
Xbit_r92_c53 bl_53 br_53 wl_92 vdd gnd cell_6t
Xbit_r93_c53 bl_53 br_53 wl_93 vdd gnd cell_6t
Xbit_r94_c53 bl_53 br_53 wl_94 vdd gnd cell_6t
Xbit_r95_c53 bl_53 br_53 wl_95 vdd gnd cell_6t
Xbit_r96_c53 bl_53 br_53 wl_96 vdd gnd cell_6t
Xbit_r97_c53 bl_53 br_53 wl_97 vdd gnd cell_6t
Xbit_r98_c53 bl_53 br_53 wl_98 vdd gnd cell_6t
Xbit_r99_c53 bl_53 br_53 wl_99 vdd gnd cell_6t
Xbit_r100_c53 bl_53 br_53 wl_100 vdd gnd cell_6t
Xbit_r101_c53 bl_53 br_53 wl_101 vdd gnd cell_6t
Xbit_r102_c53 bl_53 br_53 wl_102 vdd gnd cell_6t
Xbit_r103_c53 bl_53 br_53 wl_103 vdd gnd cell_6t
Xbit_r104_c53 bl_53 br_53 wl_104 vdd gnd cell_6t
Xbit_r105_c53 bl_53 br_53 wl_105 vdd gnd cell_6t
Xbit_r106_c53 bl_53 br_53 wl_106 vdd gnd cell_6t
Xbit_r107_c53 bl_53 br_53 wl_107 vdd gnd cell_6t
Xbit_r108_c53 bl_53 br_53 wl_108 vdd gnd cell_6t
Xbit_r109_c53 bl_53 br_53 wl_109 vdd gnd cell_6t
Xbit_r110_c53 bl_53 br_53 wl_110 vdd gnd cell_6t
Xbit_r111_c53 bl_53 br_53 wl_111 vdd gnd cell_6t
Xbit_r112_c53 bl_53 br_53 wl_112 vdd gnd cell_6t
Xbit_r113_c53 bl_53 br_53 wl_113 vdd gnd cell_6t
Xbit_r114_c53 bl_53 br_53 wl_114 vdd gnd cell_6t
Xbit_r115_c53 bl_53 br_53 wl_115 vdd gnd cell_6t
Xbit_r116_c53 bl_53 br_53 wl_116 vdd gnd cell_6t
Xbit_r117_c53 bl_53 br_53 wl_117 vdd gnd cell_6t
Xbit_r118_c53 bl_53 br_53 wl_118 vdd gnd cell_6t
Xbit_r119_c53 bl_53 br_53 wl_119 vdd gnd cell_6t
Xbit_r120_c53 bl_53 br_53 wl_120 vdd gnd cell_6t
Xbit_r121_c53 bl_53 br_53 wl_121 vdd gnd cell_6t
Xbit_r122_c53 bl_53 br_53 wl_122 vdd gnd cell_6t
Xbit_r123_c53 bl_53 br_53 wl_123 vdd gnd cell_6t
Xbit_r124_c53 bl_53 br_53 wl_124 vdd gnd cell_6t
Xbit_r125_c53 bl_53 br_53 wl_125 vdd gnd cell_6t
Xbit_r126_c53 bl_53 br_53 wl_126 vdd gnd cell_6t
Xbit_r127_c53 bl_53 br_53 wl_127 vdd gnd cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd cell_6t
Xbit_r1_c54 bl_54 br_54 wl_1 vdd gnd cell_6t
Xbit_r2_c54 bl_54 br_54 wl_2 vdd gnd cell_6t
Xbit_r3_c54 bl_54 br_54 wl_3 vdd gnd cell_6t
Xbit_r4_c54 bl_54 br_54 wl_4 vdd gnd cell_6t
Xbit_r5_c54 bl_54 br_54 wl_5 vdd gnd cell_6t
Xbit_r6_c54 bl_54 br_54 wl_6 vdd gnd cell_6t
Xbit_r7_c54 bl_54 br_54 wl_7 vdd gnd cell_6t
Xbit_r8_c54 bl_54 br_54 wl_8 vdd gnd cell_6t
Xbit_r9_c54 bl_54 br_54 wl_9 vdd gnd cell_6t
Xbit_r10_c54 bl_54 br_54 wl_10 vdd gnd cell_6t
Xbit_r11_c54 bl_54 br_54 wl_11 vdd gnd cell_6t
Xbit_r12_c54 bl_54 br_54 wl_12 vdd gnd cell_6t
Xbit_r13_c54 bl_54 br_54 wl_13 vdd gnd cell_6t
Xbit_r14_c54 bl_54 br_54 wl_14 vdd gnd cell_6t
Xbit_r15_c54 bl_54 br_54 wl_15 vdd gnd cell_6t
Xbit_r16_c54 bl_54 br_54 wl_16 vdd gnd cell_6t
Xbit_r17_c54 bl_54 br_54 wl_17 vdd gnd cell_6t
Xbit_r18_c54 bl_54 br_54 wl_18 vdd gnd cell_6t
Xbit_r19_c54 bl_54 br_54 wl_19 vdd gnd cell_6t
Xbit_r20_c54 bl_54 br_54 wl_20 vdd gnd cell_6t
Xbit_r21_c54 bl_54 br_54 wl_21 vdd gnd cell_6t
Xbit_r22_c54 bl_54 br_54 wl_22 vdd gnd cell_6t
Xbit_r23_c54 bl_54 br_54 wl_23 vdd gnd cell_6t
Xbit_r24_c54 bl_54 br_54 wl_24 vdd gnd cell_6t
Xbit_r25_c54 bl_54 br_54 wl_25 vdd gnd cell_6t
Xbit_r26_c54 bl_54 br_54 wl_26 vdd gnd cell_6t
Xbit_r27_c54 bl_54 br_54 wl_27 vdd gnd cell_6t
Xbit_r28_c54 bl_54 br_54 wl_28 vdd gnd cell_6t
Xbit_r29_c54 bl_54 br_54 wl_29 vdd gnd cell_6t
Xbit_r30_c54 bl_54 br_54 wl_30 vdd gnd cell_6t
Xbit_r31_c54 bl_54 br_54 wl_31 vdd gnd cell_6t
Xbit_r32_c54 bl_54 br_54 wl_32 vdd gnd cell_6t
Xbit_r33_c54 bl_54 br_54 wl_33 vdd gnd cell_6t
Xbit_r34_c54 bl_54 br_54 wl_34 vdd gnd cell_6t
Xbit_r35_c54 bl_54 br_54 wl_35 vdd gnd cell_6t
Xbit_r36_c54 bl_54 br_54 wl_36 vdd gnd cell_6t
Xbit_r37_c54 bl_54 br_54 wl_37 vdd gnd cell_6t
Xbit_r38_c54 bl_54 br_54 wl_38 vdd gnd cell_6t
Xbit_r39_c54 bl_54 br_54 wl_39 vdd gnd cell_6t
Xbit_r40_c54 bl_54 br_54 wl_40 vdd gnd cell_6t
Xbit_r41_c54 bl_54 br_54 wl_41 vdd gnd cell_6t
Xbit_r42_c54 bl_54 br_54 wl_42 vdd gnd cell_6t
Xbit_r43_c54 bl_54 br_54 wl_43 vdd gnd cell_6t
Xbit_r44_c54 bl_54 br_54 wl_44 vdd gnd cell_6t
Xbit_r45_c54 bl_54 br_54 wl_45 vdd gnd cell_6t
Xbit_r46_c54 bl_54 br_54 wl_46 vdd gnd cell_6t
Xbit_r47_c54 bl_54 br_54 wl_47 vdd gnd cell_6t
Xbit_r48_c54 bl_54 br_54 wl_48 vdd gnd cell_6t
Xbit_r49_c54 bl_54 br_54 wl_49 vdd gnd cell_6t
Xbit_r50_c54 bl_54 br_54 wl_50 vdd gnd cell_6t
Xbit_r51_c54 bl_54 br_54 wl_51 vdd gnd cell_6t
Xbit_r52_c54 bl_54 br_54 wl_52 vdd gnd cell_6t
Xbit_r53_c54 bl_54 br_54 wl_53 vdd gnd cell_6t
Xbit_r54_c54 bl_54 br_54 wl_54 vdd gnd cell_6t
Xbit_r55_c54 bl_54 br_54 wl_55 vdd gnd cell_6t
Xbit_r56_c54 bl_54 br_54 wl_56 vdd gnd cell_6t
Xbit_r57_c54 bl_54 br_54 wl_57 vdd gnd cell_6t
Xbit_r58_c54 bl_54 br_54 wl_58 vdd gnd cell_6t
Xbit_r59_c54 bl_54 br_54 wl_59 vdd gnd cell_6t
Xbit_r60_c54 bl_54 br_54 wl_60 vdd gnd cell_6t
Xbit_r61_c54 bl_54 br_54 wl_61 vdd gnd cell_6t
Xbit_r62_c54 bl_54 br_54 wl_62 vdd gnd cell_6t
Xbit_r63_c54 bl_54 br_54 wl_63 vdd gnd cell_6t
Xbit_r64_c54 bl_54 br_54 wl_64 vdd gnd cell_6t
Xbit_r65_c54 bl_54 br_54 wl_65 vdd gnd cell_6t
Xbit_r66_c54 bl_54 br_54 wl_66 vdd gnd cell_6t
Xbit_r67_c54 bl_54 br_54 wl_67 vdd gnd cell_6t
Xbit_r68_c54 bl_54 br_54 wl_68 vdd gnd cell_6t
Xbit_r69_c54 bl_54 br_54 wl_69 vdd gnd cell_6t
Xbit_r70_c54 bl_54 br_54 wl_70 vdd gnd cell_6t
Xbit_r71_c54 bl_54 br_54 wl_71 vdd gnd cell_6t
Xbit_r72_c54 bl_54 br_54 wl_72 vdd gnd cell_6t
Xbit_r73_c54 bl_54 br_54 wl_73 vdd gnd cell_6t
Xbit_r74_c54 bl_54 br_54 wl_74 vdd gnd cell_6t
Xbit_r75_c54 bl_54 br_54 wl_75 vdd gnd cell_6t
Xbit_r76_c54 bl_54 br_54 wl_76 vdd gnd cell_6t
Xbit_r77_c54 bl_54 br_54 wl_77 vdd gnd cell_6t
Xbit_r78_c54 bl_54 br_54 wl_78 vdd gnd cell_6t
Xbit_r79_c54 bl_54 br_54 wl_79 vdd gnd cell_6t
Xbit_r80_c54 bl_54 br_54 wl_80 vdd gnd cell_6t
Xbit_r81_c54 bl_54 br_54 wl_81 vdd gnd cell_6t
Xbit_r82_c54 bl_54 br_54 wl_82 vdd gnd cell_6t
Xbit_r83_c54 bl_54 br_54 wl_83 vdd gnd cell_6t
Xbit_r84_c54 bl_54 br_54 wl_84 vdd gnd cell_6t
Xbit_r85_c54 bl_54 br_54 wl_85 vdd gnd cell_6t
Xbit_r86_c54 bl_54 br_54 wl_86 vdd gnd cell_6t
Xbit_r87_c54 bl_54 br_54 wl_87 vdd gnd cell_6t
Xbit_r88_c54 bl_54 br_54 wl_88 vdd gnd cell_6t
Xbit_r89_c54 bl_54 br_54 wl_89 vdd gnd cell_6t
Xbit_r90_c54 bl_54 br_54 wl_90 vdd gnd cell_6t
Xbit_r91_c54 bl_54 br_54 wl_91 vdd gnd cell_6t
Xbit_r92_c54 bl_54 br_54 wl_92 vdd gnd cell_6t
Xbit_r93_c54 bl_54 br_54 wl_93 vdd gnd cell_6t
Xbit_r94_c54 bl_54 br_54 wl_94 vdd gnd cell_6t
Xbit_r95_c54 bl_54 br_54 wl_95 vdd gnd cell_6t
Xbit_r96_c54 bl_54 br_54 wl_96 vdd gnd cell_6t
Xbit_r97_c54 bl_54 br_54 wl_97 vdd gnd cell_6t
Xbit_r98_c54 bl_54 br_54 wl_98 vdd gnd cell_6t
Xbit_r99_c54 bl_54 br_54 wl_99 vdd gnd cell_6t
Xbit_r100_c54 bl_54 br_54 wl_100 vdd gnd cell_6t
Xbit_r101_c54 bl_54 br_54 wl_101 vdd gnd cell_6t
Xbit_r102_c54 bl_54 br_54 wl_102 vdd gnd cell_6t
Xbit_r103_c54 bl_54 br_54 wl_103 vdd gnd cell_6t
Xbit_r104_c54 bl_54 br_54 wl_104 vdd gnd cell_6t
Xbit_r105_c54 bl_54 br_54 wl_105 vdd gnd cell_6t
Xbit_r106_c54 bl_54 br_54 wl_106 vdd gnd cell_6t
Xbit_r107_c54 bl_54 br_54 wl_107 vdd gnd cell_6t
Xbit_r108_c54 bl_54 br_54 wl_108 vdd gnd cell_6t
Xbit_r109_c54 bl_54 br_54 wl_109 vdd gnd cell_6t
Xbit_r110_c54 bl_54 br_54 wl_110 vdd gnd cell_6t
Xbit_r111_c54 bl_54 br_54 wl_111 vdd gnd cell_6t
Xbit_r112_c54 bl_54 br_54 wl_112 vdd gnd cell_6t
Xbit_r113_c54 bl_54 br_54 wl_113 vdd gnd cell_6t
Xbit_r114_c54 bl_54 br_54 wl_114 vdd gnd cell_6t
Xbit_r115_c54 bl_54 br_54 wl_115 vdd gnd cell_6t
Xbit_r116_c54 bl_54 br_54 wl_116 vdd gnd cell_6t
Xbit_r117_c54 bl_54 br_54 wl_117 vdd gnd cell_6t
Xbit_r118_c54 bl_54 br_54 wl_118 vdd gnd cell_6t
Xbit_r119_c54 bl_54 br_54 wl_119 vdd gnd cell_6t
Xbit_r120_c54 bl_54 br_54 wl_120 vdd gnd cell_6t
Xbit_r121_c54 bl_54 br_54 wl_121 vdd gnd cell_6t
Xbit_r122_c54 bl_54 br_54 wl_122 vdd gnd cell_6t
Xbit_r123_c54 bl_54 br_54 wl_123 vdd gnd cell_6t
Xbit_r124_c54 bl_54 br_54 wl_124 vdd gnd cell_6t
Xbit_r125_c54 bl_54 br_54 wl_125 vdd gnd cell_6t
Xbit_r126_c54 bl_54 br_54 wl_126 vdd gnd cell_6t
Xbit_r127_c54 bl_54 br_54 wl_127 vdd gnd cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd cell_6t
Xbit_r1_c55 bl_55 br_55 wl_1 vdd gnd cell_6t
Xbit_r2_c55 bl_55 br_55 wl_2 vdd gnd cell_6t
Xbit_r3_c55 bl_55 br_55 wl_3 vdd gnd cell_6t
Xbit_r4_c55 bl_55 br_55 wl_4 vdd gnd cell_6t
Xbit_r5_c55 bl_55 br_55 wl_5 vdd gnd cell_6t
Xbit_r6_c55 bl_55 br_55 wl_6 vdd gnd cell_6t
Xbit_r7_c55 bl_55 br_55 wl_7 vdd gnd cell_6t
Xbit_r8_c55 bl_55 br_55 wl_8 vdd gnd cell_6t
Xbit_r9_c55 bl_55 br_55 wl_9 vdd gnd cell_6t
Xbit_r10_c55 bl_55 br_55 wl_10 vdd gnd cell_6t
Xbit_r11_c55 bl_55 br_55 wl_11 vdd gnd cell_6t
Xbit_r12_c55 bl_55 br_55 wl_12 vdd gnd cell_6t
Xbit_r13_c55 bl_55 br_55 wl_13 vdd gnd cell_6t
Xbit_r14_c55 bl_55 br_55 wl_14 vdd gnd cell_6t
Xbit_r15_c55 bl_55 br_55 wl_15 vdd gnd cell_6t
Xbit_r16_c55 bl_55 br_55 wl_16 vdd gnd cell_6t
Xbit_r17_c55 bl_55 br_55 wl_17 vdd gnd cell_6t
Xbit_r18_c55 bl_55 br_55 wl_18 vdd gnd cell_6t
Xbit_r19_c55 bl_55 br_55 wl_19 vdd gnd cell_6t
Xbit_r20_c55 bl_55 br_55 wl_20 vdd gnd cell_6t
Xbit_r21_c55 bl_55 br_55 wl_21 vdd gnd cell_6t
Xbit_r22_c55 bl_55 br_55 wl_22 vdd gnd cell_6t
Xbit_r23_c55 bl_55 br_55 wl_23 vdd gnd cell_6t
Xbit_r24_c55 bl_55 br_55 wl_24 vdd gnd cell_6t
Xbit_r25_c55 bl_55 br_55 wl_25 vdd gnd cell_6t
Xbit_r26_c55 bl_55 br_55 wl_26 vdd gnd cell_6t
Xbit_r27_c55 bl_55 br_55 wl_27 vdd gnd cell_6t
Xbit_r28_c55 bl_55 br_55 wl_28 vdd gnd cell_6t
Xbit_r29_c55 bl_55 br_55 wl_29 vdd gnd cell_6t
Xbit_r30_c55 bl_55 br_55 wl_30 vdd gnd cell_6t
Xbit_r31_c55 bl_55 br_55 wl_31 vdd gnd cell_6t
Xbit_r32_c55 bl_55 br_55 wl_32 vdd gnd cell_6t
Xbit_r33_c55 bl_55 br_55 wl_33 vdd gnd cell_6t
Xbit_r34_c55 bl_55 br_55 wl_34 vdd gnd cell_6t
Xbit_r35_c55 bl_55 br_55 wl_35 vdd gnd cell_6t
Xbit_r36_c55 bl_55 br_55 wl_36 vdd gnd cell_6t
Xbit_r37_c55 bl_55 br_55 wl_37 vdd gnd cell_6t
Xbit_r38_c55 bl_55 br_55 wl_38 vdd gnd cell_6t
Xbit_r39_c55 bl_55 br_55 wl_39 vdd gnd cell_6t
Xbit_r40_c55 bl_55 br_55 wl_40 vdd gnd cell_6t
Xbit_r41_c55 bl_55 br_55 wl_41 vdd gnd cell_6t
Xbit_r42_c55 bl_55 br_55 wl_42 vdd gnd cell_6t
Xbit_r43_c55 bl_55 br_55 wl_43 vdd gnd cell_6t
Xbit_r44_c55 bl_55 br_55 wl_44 vdd gnd cell_6t
Xbit_r45_c55 bl_55 br_55 wl_45 vdd gnd cell_6t
Xbit_r46_c55 bl_55 br_55 wl_46 vdd gnd cell_6t
Xbit_r47_c55 bl_55 br_55 wl_47 vdd gnd cell_6t
Xbit_r48_c55 bl_55 br_55 wl_48 vdd gnd cell_6t
Xbit_r49_c55 bl_55 br_55 wl_49 vdd gnd cell_6t
Xbit_r50_c55 bl_55 br_55 wl_50 vdd gnd cell_6t
Xbit_r51_c55 bl_55 br_55 wl_51 vdd gnd cell_6t
Xbit_r52_c55 bl_55 br_55 wl_52 vdd gnd cell_6t
Xbit_r53_c55 bl_55 br_55 wl_53 vdd gnd cell_6t
Xbit_r54_c55 bl_55 br_55 wl_54 vdd gnd cell_6t
Xbit_r55_c55 bl_55 br_55 wl_55 vdd gnd cell_6t
Xbit_r56_c55 bl_55 br_55 wl_56 vdd gnd cell_6t
Xbit_r57_c55 bl_55 br_55 wl_57 vdd gnd cell_6t
Xbit_r58_c55 bl_55 br_55 wl_58 vdd gnd cell_6t
Xbit_r59_c55 bl_55 br_55 wl_59 vdd gnd cell_6t
Xbit_r60_c55 bl_55 br_55 wl_60 vdd gnd cell_6t
Xbit_r61_c55 bl_55 br_55 wl_61 vdd gnd cell_6t
Xbit_r62_c55 bl_55 br_55 wl_62 vdd gnd cell_6t
Xbit_r63_c55 bl_55 br_55 wl_63 vdd gnd cell_6t
Xbit_r64_c55 bl_55 br_55 wl_64 vdd gnd cell_6t
Xbit_r65_c55 bl_55 br_55 wl_65 vdd gnd cell_6t
Xbit_r66_c55 bl_55 br_55 wl_66 vdd gnd cell_6t
Xbit_r67_c55 bl_55 br_55 wl_67 vdd gnd cell_6t
Xbit_r68_c55 bl_55 br_55 wl_68 vdd gnd cell_6t
Xbit_r69_c55 bl_55 br_55 wl_69 vdd gnd cell_6t
Xbit_r70_c55 bl_55 br_55 wl_70 vdd gnd cell_6t
Xbit_r71_c55 bl_55 br_55 wl_71 vdd gnd cell_6t
Xbit_r72_c55 bl_55 br_55 wl_72 vdd gnd cell_6t
Xbit_r73_c55 bl_55 br_55 wl_73 vdd gnd cell_6t
Xbit_r74_c55 bl_55 br_55 wl_74 vdd gnd cell_6t
Xbit_r75_c55 bl_55 br_55 wl_75 vdd gnd cell_6t
Xbit_r76_c55 bl_55 br_55 wl_76 vdd gnd cell_6t
Xbit_r77_c55 bl_55 br_55 wl_77 vdd gnd cell_6t
Xbit_r78_c55 bl_55 br_55 wl_78 vdd gnd cell_6t
Xbit_r79_c55 bl_55 br_55 wl_79 vdd gnd cell_6t
Xbit_r80_c55 bl_55 br_55 wl_80 vdd gnd cell_6t
Xbit_r81_c55 bl_55 br_55 wl_81 vdd gnd cell_6t
Xbit_r82_c55 bl_55 br_55 wl_82 vdd gnd cell_6t
Xbit_r83_c55 bl_55 br_55 wl_83 vdd gnd cell_6t
Xbit_r84_c55 bl_55 br_55 wl_84 vdd gnd cell_6t
Xbit_r85_c55 bl_55 br_55 wl_85 vdd gnd cell_6t
Xbit_r86_c55 bl_55 br_55 wl_86 vdd gnd cell_6t
Xbit_r87_c55 bl_55 br_55 wl_87 vdd gnd cell_6t
Xbit_r88_c55 bl_55 br_55 wl_88 vdd gnd cell_6t
Xbit_r89_c55 bl_55 br_55 wl_89 vdd gnd cell_6t
Xbit_r90_c55 bl_55 br_55 wl_90 vdd gnd cell_6t
Xbit_r91_c55 bl_55 br_55 wl_91 vdd gnd cell_6t
Xbit_r92_c55 bl_55 br_55 wl_92 vdd gnd cell_6t
Xbit_r93_c55 bl_55 br_55 wl_93 vdd gnd cell_6t
Xbit_r94_c55 bl_55 br_55 wl_94 vdd gnd cell_6t
Xbit_r95_c55 bl_55 br_55 wl_95 vdd gnd cell_6t
Xbit_r96_c55 bl_55 br_55 wl_96 vdd gnd cell_6t
Xbit_r97_c55 bl_55 br_55 wl_97 vdd gnd cell_6t
Xbit_r98_c55 bl_55 br_55 wl_98 vdd gnd cell_6t
Xbit_r99_c55 bl_55 br_55 wl_99 vdd gnd cell_6t
Xbit_r100_c55 bl_55 br_55 wl_100 vdd gnd cell_6t
Xbit_r101_c55 bl_55 br_55 wl_101 vdd gnd cell_6t
Xbit_r102_c55 bl_55 br_55 wl_102 vdd gnd cell_6t
Xbit_r103_c55 bl_55 br_55 wl_103 vdd gnd cell_6t
Xbit_r104_c55 bl_55 br_55 wl_104 vdd gnd cell_6t
Xbit_r105_c55 bl_55 br_55 wl_105 vdd gnd cell_6t
Xbit_r106_c55 bl_55 br_55 wl_106 vdd gnd cell_6t
Xbit_r107_c55 bl_55 br_55 wl_107 vdd gnd cell_6t
Xbit_r108_c55 bl_55 br_55 wl_108 vdd gnd cell_6t
Xbit_r109_c55 bl_55 br_55 wl_109 vdd gnd cell_6t
Xbit_r110_c55 bl_55 br_55 wl_110 vdd gnd cell_6t
Xbit_r111_c55 bl_55 br_55 wl_111 vdd gnd cell_6t
Xbit_r112_c55 bl_55 br_55 wl_112 vdd gnd cell_6t
Xbit_r113_c55 bl_55 br_55 wl_113 vdd gnd cell_6t
Xbit_r114_c55 bl_55 br_55 wl_114 vdd gnd cell_6t
Xbit_r115_c55 bl_55 br_55 wl_115 vdd gnd cell_6t
Xbit_r116_c55 bl_55 br_55 wl_116 vdd gnd cell_6t
Xbit_r117_c55 bl_55 br_55 wl_117 vdd gnd cell_6t
Xbit_r118_c55 bl_55 br_55 wl_118 vdd gnd cell_6t
Xbit_r119_c55 bl_55 br_55 wl_119 vdd gnd cell_6t
Xbit_r120_c55 bl_55 br_55 wl_120 vdd gnd cell_6t
Xbit_r121_c55 bl_55 br_55 wl_121 vdd gnd cell_6t
Xbit_r122_c55 bl_55 br_55 wl_122 vdd gnd cell_6t
Xbit_r123_c55 bl_55 br_55 wl_123 vdd gnd cell_6t
Xbit_r124_c55 bl_55 br_55 wl_124 vdd gnd cell_6t
Xbit_r125_c55 bl_55 br_55 wl_125 vdd gnd cell_6t
Xbit_r126_c55 bl_55 br_55 wl_126 vdd gnd cell_6t
Xbit_r127_c55 bl_55 br_55 wl_127 vdd gnd cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd cell_6t
Xbit_r1_c56 bl_56 br_56 wl_1 vdd gnd cell_6t
Xbit_r2_c56 bl_56 br_56 wl_2 vdd gnd cell_6t
Xbit_r3_c56 bl_56 br_56 wl_3 vdd gnd cell_6t
Xbit_r4_c56 bl_56 br_56 wl_4 vdd gnd cell_6t
Xbit_r5_c56 bl_56 br_56 wl_5 vdd gnd cell_6t
Xbit_r6_c56 bl_56 br_56 wl_6 vdd gnd cell_6t
Xbit_r7_c56 bl_56 br_56 wl_7 vdd gnd cell_6t
Xbit_r8_c56 bl_56 br_56 wl_8 vdd gnd cell_6t
Xbit_r9_c56 bl_56 br_56 wl_9 vdd gnd cell_6t
Xbit_r10_c56 bl_56 br_56 wl_10 vdd gnd cell_6t
Xbit_r11_c56 bl_56 br_56 wl_11 vdd gnd cell_6t
Xbit_r12_c56 bl_56 br_56 wl_12 vdd gnd cell_6t
Xbit_r13_c56 bl_56 br_56 wl_13 vdd gnd cell_6t
Xbit_r14_c56 bl_56 br_56 wl_14 vdd gnd cell_6t
Xbit_r15_c56 bl_56 br_56 wl_15 vdd gnd cell_6t
Xbit_r16_c56 bl_56 br_56 wl_16 vdd gnd cell_6t
Xbit_r17_c56 bl_56 br_56 wl_17 vdd gnd cell_6t
Xbit_r18_c56 bl_56 br_56 wl_18 vdd gnd cell_6t
Xbit_r19_c56 bl_56 br_56 wl_19 vdd gnd cell_6t
Xbit_r20_c56 bl_56 br_56 wl_20 vdd gnd cell_6t
Xbit_r21_c56 bl_56 br_56 wl_21 vdd gnd cell_6t
Xbit_r22_c56 bl_56 br_56 wl_22 vdd gnd cell_6t
Xbit_r23_c56 bl_56 br_56 wl_23 vdd gnd cell_6t
Xbit_r24_c56 bl_56 br_56 wl_24 vdd gnd cell_6t
Xbit_r25_c56 bl_56 br_56 wl_25 vdd gnd cell_6t
Xbit_r26_c56 bl_56 br_56 wl_26 vdd gnd cell_6t
Xbit_r27_c56 bl_56 br_56 wl_27 vdd gnd cell_6t
Xbit_r28_c56 bl_56 br_56 wl_28 vdd gnd cell_6t
Xbit_r29_c56 bl_56 br_56 wl_29 vdd gnd cell_6t
Xbit_r30_c56 bl_56 br_56 wl_30 vdd gnd cell_6t
Xbit_r31_c56 bl_56 br_56 wl_31 vdd gnd cell_6t
Xbit_r32_c56 bl_56 br_56 wl_32 vdd gnd cell_6t
Xbit_r33_c56 bl_56 br_56 wl_33 vdd gnd cell_6t
Xbit_r34_c56 bl_56 br_56 wl_34 vdd gnd cell_6t
Xbit_r35_c56 bl_56 br_56 wl_35 vdd gnd cell_6t
Xbit_r36_c56 bl_56 br_56 wl_36 vdd gnd cell_6t
Xbit_r37_c56 bl_56 br_56 wl_37 vdd gnd cell_6t
Xbit_r38_c56 bl_56 br_56 wl_38 vdd gnd cell_6t
Xbit_r39_c56 bl_56 br_56 wl_39 vdd gnd cell_6t
Xbit_r40_c56 bl_56 br_56 wl_40 vdd gnd cell_6t
Xbit_r41_c56 bl_56 br_56 wl_41 vdd gnd cell_6t
Xbit_r42_c56 bl_56 br_56 wl_42 vdd gnd cell_6t
Xbit_r43_c56 bl_56 br_56 wl_43 vdd gnd cell_6t
Xbit_r44_c56 bl_56 br_56 wl_44 vdd gnd cell_6t
Xbit_r45_c56 bl_56 br_56 wl_45 vdd gnd cell_6t
Xbit_r46_c56 bl_56 br_56 wl_46 vdd gnd cell_6t
Xbit_r47_c56 bl_56 br_56 wl_47 vdd gnd cell_6t
Xbit_r48_c56 bl_56 br_56 wl_48 vdd gnd cell_6t
Xbit_r49_c56 bl_56 br_56 wl_49 vdd gnd cell_6t
Xbit_r50_c56 bl_56 br_56 wl_50 vdd gnd cell_6t
Xbit_r51_c56 bl_56 br_56 wl_51 vdd gnd cell_6t
Xbit_r52_c56 bl_56 br_56 wl_52 vdd gnd cell_6t
Xbit_r53_c56 bl_56 br_56 wl_53 vdd gnd cell_6t
Xbit_r54_c56 bl_56 br_56 wl_54 vdd gnd cell_6t
Xbit_r55_c56 bl_56 br_56 wl_55 vdd gnd cell_6t
Xbit_r56_c56 bl_56 br_56 wl_56 vdd gnd cell_6t
Xbit_r57_c56 bl_56 br_56 wl_57 vdd gnd cell_6t
Xbit_r58_c56 bl_56 br_56 wl_58 vdd gnd cell_6t
Xbit_r59_c56 bl_56 br_56 wl_59 vdd gnd cell_6t
Xbit_r60_c56 bl_56 br_56 wl_60 vdd gnd cell_6t
Xbit_r61_c56 bl_56 br_56 wl_61 vdd gnd cell_6t
Xbit_r62_c56 bl_56 br_56 wl_62 vdd gnd cell_6t
Xbit_r63_c56 bl_56 br_56 wl_63 vdd gnd cell_6t
Xbit_r64_c56 bl_56 br_56 wl_64 vdd gnd cell_6t
Xbit_r65_c56 bl_56 br_56 wl_65 vdd gnd cell_6t
Xbit_r66_c56 bl_56 br_56 wl_66 vdd gnd cell_6t
Xbit_r67_c56 bl_56 br_56 wl_67 vdd gnd cell_6t
Xbit_r68_c56 bl_56 br_56 wl_68 vdd gnd cell_6t
Xbit_r69_c56 bl_56 br_56 wl_69 vdd gnd cell_6t
Xbit_r70_c56 bl_56 br_56 wl_70 vdd gnd cell_6t
Xbit_r71_c56 bl_56 br_56 wl_71 vdd gnd cell_6t
Xbit_r72_c56 bl_56 br_56 wl_72 vdd gnd cell_6t
Xbit_r73_c56 bl_56 br_56 wl_73 vdd gnd cell_6t
Xbit_r74_c56 bl_56 br_56 wl_74 vdd gnd cell_6t
Xbit_r75_c56 bl_56 br_56 wl_75 vdd gnd cell_6t
Xbit_r76_c56 bl_56 br_56 wl_76 vdd gnd cell_6t
Xbit_r77_c56 bl_56 br_56 wl_77 vdd gnd cell_6t
Xbit_r78_c56 bl_56 br_56 wl_78 vdd gnd cell_6t
Xbit_r79_c56 bl_56 br_56 wl_79 vdd gnd cell_6t
Xbit_r80_c56 bl_56 br_56 wl_80 vdd gnd cell_6t
Xbit_r81_c56 bl_56 br_56 wl_81 vdd gnd cell_6t
Xbit_r82_c56 bl_56 br_56 wl_82 vdd gnd cell_6t
Xbit_r83_c56 bl_56 br_56 wl_83 vdd gnd cell_6t
Xbit_r84_c56 bl_56 br_56 wl_84 vdd gnd cell_6t
Xbit_r85_c56 bl_56 br_56 wl_85 vdd gnd cell_6t
Xbit_r86_c56 bl_56 br_56 wl_86 vdd gnd cell_6t
Xbit_r87_c56 bl_56 br_56 wl_87 vdd gnd cell_6t
Xbit_r88_c56 bl_56 br_56 wl_88 vdd gnd cell_6t
Xbit_r89_c56 bl_56 br_56 wl_89 vdd gnd cell_6t
Xbit_r90_c56 bl_56 br_56 wl_90 vdd gnd cell_6t
Xbit_r91_c56 bl_56 br_56 wl_91 vdd gnd cell_6t
Xbit_r92_c56 bl_56 br_56 wl_92 vdd gnd cell_6t
Xbit_r93_c56 bl_56 br_56 wl_93 vdd gnd cell_6t
Xbit_r94_c56 bl_56 br_56 wl_94 vdd gnd cell_6t
Xbit_r95_c56 bl_56 br_56 wl_95 vdd gnd cell_6t
Xbit_r96_c56 bl_56 br_56 wl_96 vdd gnd cell_6t
Xbit_r97_c56 bl_56 br_56 wl_97 vdd gnd cell_6t
Xbit_r98_c56 bl_56 br_56 wl_98 vdd gnd cell_6t
Xbit_r99_c56 bl_56 br_56 wl_99 vdd gnd cell_6t
Xbit_r100_c56 bl_56 br_56 wl_100 vdd gnd cell_6t
Xbit_r101_c56 bl_56 br_56 wl_101 vdd gnd cell_6t
Xbit_r102_c56 bl_56 br_56 wl_102 vdd gnd cell_6t
Xbit_r103_c56 bl_56 br_56 wl_103 vdd gnd cell_6t
Xbit_r104_c56 bl_56 br_56 wl_104 vdd gnd cell_6t
Xbit_r105_c56 bl_56 br_56 wl_105 vdd gnd cell_6t
Xbit_r106_c56 bl_56 br_56 wl_106 vdd gnd cell_6t
Xbit_r107_c56 bl_56 br_56 wl_107 vdd gnd cell_6t
Xbit_r108_c56 bl_56 br_56 wl_108 vdd gnd cell_6t
Xbit_r109_c56 bl_56 br_56 wl_109 vdd gnd cell_6t
Xbit_r110_c56 bl_56 br_56 wl_110 vdd gnd cell_6t
Xbit_r111_c56 bl_56 br_56 wl_111 vdd gnd cell_6t
Xbit_r112_c56 bl_56 br_56 wl_112 vdd gnd cell_6t
Xbit_r113_c56 bl_56 br_56 wl_113 vdd gnd cell_6t
Xbit_r114_c56 bl_56 br_56 wl_114 vdd gnd cell_6t
Xbit_r115_c56 bl_56 br_56 wl_115 vdd gnd cell_6t
Xbit_r116_c56 bl_56 br_56 wl_116 vdd gnd cell_6t
Xbit_r117_c56 bl_56 br_56 wl_117 vdd gnd cell_6t
Xbit_r118_c56 bl_56 br_56 wl_118 vdd gnd cell_6t
Xbit_r119_c56 bl_56 br_56 wl_119 vdd gnd cell_6t
Xbit_r120_c56 bl_56 br_56 wl_120 vdd gnd cell_6t
Xbit_r121_c56 bl_56 br_56 wl_121 vdd gnd cell_6t
Xbit_r122_c56 bl_56 br_56 wl_122 vdd gnd cell_6t
Xbit_r123_c56 bl_56 br_56 wl_123 vdd gnd cell_6t
Xbit_r124_c56 bl_56 br_56 wl_124 vdd gnd cell_6t
Xbit_r125_c56 bl_56 br_56 wl_125 vdd gnd cell_6t
Xbit_r126_c56 bl_56 br_56 wl_126 vdd gnd cell_6t
Xbit_r127_c56 bl_56 br_56 wl_127 vdd gnd cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd cell_6t
Xbit_r1_c57 bl_57 br_57 wl_1 vdd gnd cell_6t
Xbit_r2_c57 bl_57 br_57 wl_2 vdd gnd cell_6t
Xbit_r3_c57 bl_57 br_57 wl_3 vdd gnd cell_6t
Xbit_r4_c57 bl_57 br_57 wl_4 vdd gnd cell_6t
Xbit_r5_c57 bl_57 br_57 wl_5 vdd gnd cell_6t
Xbit_r6_c57 bl_57 br_57 wl_6 vdd gnd cell_6t
Xbit_r7_c57 bl_57 br_57 wl_7 vdd gnd cell_6t
Xbit_r8_c57 bl_57 br_57 wl_8 vdd gnd cell_6t
Xbit_r9_c57 bl_57 br_57 wl_9 vdd gnd cell_6t
Xbit_r10_c57 bl_57 br_57 wl_10 vdd gnd cell_6t
Xbit_r11_c57 bl_57 br_57 wl_11 vdd gnd cell_6t
Xbit_r12_c57 bl_57 br_57 wl_12 vdd gnd cell_6t
Xbit_r13_c57 bl_57 br_57 wl_13 vdd gnd cell_6t
Xbit_r14_c57 bl_57 br_57 wl_14 vdd gnd cell_6t
Xbit_r15_c57 bl_57 br_57 wl_15 vdd gnd cell_6t
Xbit_r16_c57 bl_57 br_57 wl_16 vdd gnd cell_6t
Xbit_r17_c57 bl_57 br_57 wl_17 vdd gnd cell_6t
Xbit_r18_c57 bl_57 br_57 wl_18 vdd gnd cell_6t
Xbit_r19_c57 bl_57 br_57 wl_19 vdd gnd cell_6t
Xbit_r20_c57 bl_57 br_57 wl_20 vdd gnd cell_6t
Xbit_r21_c57 bl_57 br_57 wl_21 vdd gnd cell_6t
Xbit_r22_c57 bl_57 br_57 wl_22 vdd gnd cell_6t
Xbit_r23_c57 bl_57 br_57 wl_23 vdd gnd cell_6t
Xbit_r24_c57 bl_57 br_57 wl_24 vdd gnd cell_6t
Xbit_r25_c57 bl_57 br_57 wl_25 vdd gnd cell_6t
Xbit_r26_c57 bl_57 br_57 wl_26 vdd gnd cell_6t
Xbit_r27_c57 bl_57 br_57 wl_27 vdd gnd cell_6t
Xbit_r28_c57 bl_57 br_57 wl_28 vdd gnd cell_6t
Xbit_r29_c57 bl_57 br_57 wl_29 vdd gnd cell_6t
Xbit_r30_c57 bl_57 br_57 wl_30 vdd gnd cell_6t
Xbit_r31_c57 bl_57 br_57 wl_31 vdd gnd cell_6t
Xbit_r32_c57 bl_57 br_57 wl_32 vdd gnd cell_6t
Xbit_r33_c57 bl_57 br_57 wl_33 vdd gnd cell_6t
Xbit_r34_c57 bl_57 br_57 wl_34 vdd gnd cell_6t
Xbit_r35_c57 bl_57 br_57 wl_35 vdd gnd cell_6t
Xbit_r36_c57 bl_57 br_57 wl_36 vdd gnd cell_6t
Xbit_r37_c57 bl_57 br_57 wl_37 vdd gnd cell_6t
Xbit_r38_c57 bl_57 br_57 wl_38 vdd gnd cell_6t
Xbit_r39_c57 bl_57 br_57 wl_39 vdd gnd cell_6t
Xbit_r40_c57 bl_57 br_57 wl_40 vdd gnd cell_6t
Xbit_r41_c57 bl_57 br_57 wl_41 vdd gnd cell_6t
Xbit_r42_c57 bl_57 br_57 wl_42 vdd gnd cell_6t
Xbit_r43_c57 bl_57 br_57 wl_43 vdd gnd cell_6t
Xbit_r44_c57 bl_57 br_57 wl_44 vdd gnd cell_6t
Xbit_r45_c57 bl_57 br_57 wl_45 vdd gnd cell_6t
Xbit_r46_c57 bl_57 br_57 wl_46 vdd gnd cell_6t
Xbit_r47_c57 bl_57 br_57 wl_47 vdd gnd cell_6t
Xbit_r48_c57 bl_57 br_57 wl_48 vdd gnd cell_6t
Xbit_r49_c57 bl_57 br_57 wl_49 vdd gnd cell_6t
Xbit_r50_c57 bl_57 br_57 wl_50 vdd gnd cell_6t
Xbit_r51_c57 bl_57 br_57 wl_51 vdd gnd cell_6t
Xbit_r52_c57 bl_57 br_57 wl_52 vdd gnd cell_6t
Xbit_r53_c57 bl_57 br_57 wl_53 vdd gnd cell_6t
Xbit_r54_c57 bl_57 br_57 wl_54 vdd gnd cell_6t
Xbit_r55_c57 bl_57 br_57 wl_55 vdd gnd cell_6t
Xbit_r56_c57 bl_57 br_57 wl_56 vdd gnd cell_6t
Xbit_r57_c57 bl_57 br_57 wl_57 vdd gnd cell_6t
Xbit_r58_c57 bl_57 br_57 wl_58 vdd gnd cell_6t
Xbit_r59_c57 bl_57 br_57 wl_59 vdd gnd cell_6t
Xbit_r60_c57 bl_57 br_57 wl_60 vdd gnd cell_6t
Xbit_r61_c57 bl_57 br_57 wl_61 vdd gnd cell_6t
Xbit_r62_c57 bl_57 br_57 wl_62 vdd gnd cell_6t
Xbit_r63_c57 bl_57 br_57 wl_63 vdd gnd cell_6t
Xbit_r64_c57 bl_57 br_57 wl_64 vdd gnd cell_6t
Xbit_r65_c57 bl_57 br_57 wl_65 vdd gnd cell_6t
Xbit_r66_c57 bl_57 br_57 wl_66 vdd gnd cell_6t
Xbit_r67_c57 bl_57 br_57 wl_67 vdd gnd cell_6t
Xbit_r68_c57 bl_57 br_57 wl_68 vdd gnd cell_6t
Xbit_r69_c57 bl_57 br_57 wl_69 vdd gnd cell_6t
Xbit_r70_c57 bl_57 br_57 wl_70 vdd gnd cell_6t
Xbit_r71_c57 bl_57 br_57 wl_71 vdd gnd cell_6t
Xbit_r72_c57 bl_57 br_57 wl_72 vdd gnd cell_6t
Xbit_r73_c57 bl_57 br_57 wl_73 vdd gnd cell_6t
Xbit_r74_c57 bl_57 br_57 wl_74 vdd gnd cell_6t
Xbit_r75_c57 bl_57 br_57 wl_75 vdd gnd cell_6t
Xbit_r76_c57 bl_57 br_57 wl_76 vdd gnd cell_6t
Xbit_r77_c57 bl_57 br_57 wl_77 vdd gnd cell_6t
Xbit_r78_c57 bl_57 br_57 wl_78 vdd gnd cell_6t
Xbit_r79_c57 bl_57 br_57 wl_79 vdd gnd cell_6t
Xbit_r80_c57 bl_57 br_57 wl_80 vdd gnd cell_6t
Xbit_r81_c57 bl_57 br_57 wl_81 vdd gnd cell_6t
Xbit_r82_c57 bl_57 br_57 wl_82 vdd gnd cell_6t
Xbit_r83_c57 bl_57 br_57 wl_83 vdd gnd cell_6t
Xbit_r84_c57 bl_57 br_57 wl_84 vdd gnd cell_6t
Xbit_r85_c57 bl_57 br_57 wl_85 vdd gnd cell_6t
Xbit_r86_c57 bl_57 br_57 wl_86 vdd gnd cell_6t
Xbit_r87_c57 bl_57 br_57 wl_87 vdd gnd cell_6t
Xbit_r88_c57 bl_57 br_57 wl_88 vdd gnd cell_6t
Xbit_r89_c57 bl_57 br_57 wl_89 vdd gnd cell_6t
Xbit_r90_c57 bl_57 br_57 wl_90 vdd gnd cell_6t
Xbit_r91_c57 bl_57 br_57 wl_91 vdd gnd cell_6t
Xbit_r92_c57 bl_57 br_57 wl_92 vdd gnd cell_6t
Xbit_r93_c57 bl_57 br_57 wl_93 vdd gnd cell_6t
Xbit_r94_c57 bl_57 br_57 wl_94 vdd gnd cell_6t
Xbit_r95_c57 bl_57 br_57 wl_95 vdd gnd cell_6t
Xbit_r96_c57 bl_57 br_57 wl_96 vdd gnd cell_6t
Xbit_r97_c57 bl_57 br_57 wl_97 vdd gnd cell_6t
Xbit_r98_c57 bl_57 br_57 wl_98 vdd gnd cell_6t
Xbit_r99_c57 bl_57 br_57 wl_99 vdd gnd cell_6t
Xbit_r100_c57 bl_57 br_57 wl_100 vdd gnd cell_6t
Xbit_r101_c57 bl_57 br_57 wl_101 vdd gnd cell_6t
Xbit_r102_c57 bl_57 br_57 wl_102 vdd gnd cell_6t
Xbit_r103_c57 bl_57 br_57 wl_103 vdd gnd cell_6t
Xbit_r104_c57 bl_57 br_57 wl_104 vdd gnd cell_6t
Xbit_r105_c57 bl_57 br_57 wl_105 vdd gnd cell_6t
Xbit_r106_c57 bl_57 br_57 wl_106 vdd gnd cell_6t
Xbit_r107_c57 bl_57 br_57 wl_107 vdd gnd cell_6t
Xbit_r108_c57 bl_57 br_57 wl_108 vdd gnd cell_6t
Xbit_r109_c57 bl_57 br_57 wl_109 vdd gnd cell_6t
Xbit_r110_c57 bl_57 br_57 wl_110 vdd gnd cell_6t
Xbit_r111_c57 bl_57 br_57 wl_111 vdd gnd cell_6t
Xbit_r112_c57 bl_57 br_57 wl_112 vdd gnd cell_6t
Xbit_r113_c57 bl_57 br_57 wl_113 vdd gnd cell_6t
Xbit_r114_c57 bl_57 br_57 wl_114 vdd gnd cell_6t
Xbit_r115_c57 bl_57 br_57 wl_115 vdd gnd cell_6t
Xbit_r116_c57 bl_57 br_57 wl_116 vdd gnd cell_6t
Xbit_r117_c57 bl_57 br_57 wl_117 vdd gnd cell_6t
Xbit_r118_c57 bl_57 br_57 wl_118 vdd gnd cell_6t
Xbit_r119_c57 bl_57 br_57 wl_119 vdd gnd cell_6t
Xbit_r120_c57 bl_57 br_57 wl_120 vdd gnd cell_6t
Xbit_r121_c57 bl_57 br_57 wl_121 vdd gnd cell_6t
Xbit_r122_c57 bl_57 br_57 wl_122 vdd gnd cell_6t
Xbit_r123_c57 bl_57 br_57 wl_123 vdd gnd cell_6t
Xbit_r124_c57 bl_57 br_57 wl_124 vdd gnd cell_6t
Xbit_r125_c57 bl_57 br_57 wl_125 vdd gnd cell_6t
Xbit_r126_c57 bl_57 br_57 wl_126 vdd gnd cell_6t
Xbit_r127_c57 bl_57 br_57 wl_127 vdd gnd cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd cell_6t
Xbit_r1_c58 bl_58 br_58 wl_1 vdd gnd cell_6t
Xbit_r2_c58 bl_58 br_58 wl_2 vdd gnd cell_6t
Xbit_r3_c58 bl_58 br_58 wl_3 vdd gnd cell_6t
Xbit_r4_c58 bl_58 br_58 wl_4 vdd gnd cell_6t
Xbit_r5_c58 bl_58 br_58 wl_5 vdd gnd cell_6t
Xbit_r6_c58 bl_58 br_58 wl_6 vdd gnd cell_6t
Xbit_r7_c58 bl_58 br_58 wl_7 vdd gnd cell_6t
Xbit_r8_c58 bl_58 br_58 wl_8 vdd gnd cell_6t
Xbit_r9_c58 bl_58 br_58 wl_9 vdd gnd cell_6t
Xbit_r10_c58 bl_58 br_58 wl_10 vdd gnd cell_6t
Xbit_r11_c58 bl_58 br_58 wl_11 vdd gnd cell_6t
Xbit_r12_c58 bl_58 br_58 wl_12 vdd gnd cell_6t
Xbit_r13_c58 bl_58 br_58 wl_13 vdd gnd cell_6t
Xbit_r14_c58 bl_58 br_58 wl_14 vdd gnd cell_6t
Xbit_r15_c58 bl_58 br_58 wl_15 vdd gnd cell_6t
Xbit_r16_c58 bl_58 br_58 wl_16 vdd gnd cell_6t
Xbit_r17_c58 bl_58 br_58 wl_17 vdd gnd cell_6t
Xbit_r18_c58 bl_58 br_58 wl_18 vdd gnd cell_6t
Xbit_r19_c58 bl_58 br_58 wl_19 vdd gnd cell_6t
Xbit_r20_c58 bl_58 br_58 wl_20 vdd gnd cell_6t
Xbit_r21_c58 bl_58 br_58 wl_21 vdd gnd cell_6t
Xbit_r22_c58 bl_58 br_58 wl_22 vdd gnd cell_6t
Xbit_r23_c58 bl_58 br_58 wl_23 vdd gnd cell_6t
Xbit_r24_c58 bl_58 br_58 wl_24 vdd gnd cell_6t
Xbit_r25_c58 bl_58 br_58 wl_25 vdd gnd cell_6t
Xbit_r26_c58 bl_58 br_58 wl_26 vdd gnd cell_6t
Xbit_r27_c58 bl_58 br_58 wl_27 vdd gnd cell_6t
Xbit_r28_c58 bl_58 br_58 wl_28 vdd gnd cell_6t
Xbit_r29_c58 bl_58 br_58 wl_29 vdd gnd cell_6t
Xbit_r30_c58 bl_58 br_58 wl_30 vdd gnd cell_6t
Xbit_r31_c58 bl_58 br_58 wl_31 vdd gnd cell_6t
Xbit_r32_c58 bl_58 br_58 wl_32 vdd gnd cell_6t
Xbit_r33_c58 bl_58 br_58 wl_33 vdd gnd cell_6t
Xbit_r34_c58 bl_58 br_58 wl_34 vdd gnd cell_6t
Xbit_r35_c58 bl_58 br_58 wl_35 vdd gnd cell_6t
Xbit_r36_c58 bl_58 br_58 wl_36 vdd gnd cell_6t
Xbit_r37_c58 bl_58 br_58 wl_37 vdd gnd cell_6t
Xbit_r38_c58 bl_58 br_58 wl_38 vdd gnd cell_6t
Xbit_r39_c58 bl_58 br_58 wl_39 vdd gnd cell_6t
Xbit_r40_c58 bl_58 br_58 wl_40 vdd gnd cell_6t
Xbit_r41_c58 bl_58 br_58 wl_41 vdd gnd cell_6t
Xbit_r42_c58 bl_58 br_58 wl_42 vdd gnd cell_6t
Xbit_r43_c58 bl_58 br_58 wl_43 vdd gnd cell_6t
Xbit_r44_c58 bl_58 br_58 wl_44 vdd gnd cell_6t
Xbit_r45_c58 bl_58 br_58 wl_45 vdd gnd cell_6t
Xbit_r46_c58 bl_58 br_58 wl_46 vdd gnd cell_6t
Xbit_r47_c58 bl_58 br_58 wl_47 vdd gnd cell_6t
Xbit_r48_c58 bl_58 br_58 wl_48 vdd gnd cell_6t
Xbit_r49_c58 bl_58 br_58 wl_49 vdd gnd cell_6t
Xbit_r50_c58 bl_58 br_58 wl_50 vdd gnd cell_6t
Xbit_r51_c58 bl_58 br_58 wl_51 vdd gnd cell_6t
Xbit_r52_c58 bl_58 br_58 wl_52 vdd gnd cell_6t
Xbit_r53_c58 bl_58 br_58 wl_53 vdd gnd cell_6t
Xbit_r54_c58 bl_58 br_58 wl_54 vdd gnd cell_6t
Xbit_r55_c58 bl_58 br_58 wl_55 vdd gnd cell_6t
Xbit_r56_c58 bl_58 br_58 wl_56 vdd gnd cell_6t
Xbit_r57_c58 bl_58 br_58 wl_57 vdd gnd cell_6t
Xbit_r58_c58 bl_58 br_58 wl_58 vdd gnd cell_6t
Xbit_r59_c58 bl_58 br_58 wl_59 vdd gnd cell_6t
Xbit_r60_c58 bl_58 br_58 wl_60 vdd gnd cell_6t
Xbit_r61_c58 bl_58 br_58 wl_61 vdd gnd cell_6t
Xbit_r62_c58 bl_58 br_58 wl_62 vdd gnd cell_6t
Xbit_r63_c58 bl_58 br_58 wl_63 vdd gnd cell_6t
Xbit_r64_c58 bl_58 br_58 wl_64 vdd gnd cell_6t
Xbit_r65_c58 bl_58 br_58 wl_65 vdd gnd cell_6t
Xbit_r66_c58 bl_58 br_58 wl_66 vdd gnd cell_6t
Xbit_r67_c58 bl_58 br_58 wl_67 vdd gnd cell_6t
Xbit_r68_c58 bl_58 br_58 wl_68 vdd gnd cell_6t
Xbit_r69_c58 bl_58 br_58 wl_69 vdd gnd cell_6t
Xbit_r70_c58 bl_58 br_58 wl_70 vdd gnd cell_6t
Xbit_r71_c58 bl_58 br_58 wl_71 vdd gnd cell_6t
Xbit_r72_c58 bl_58 br_58 wl_72 vdd gnd cell_6t
Xbit_r73_c58 bl_58 br_58 wl_73 vdd gnd cell_6t
Xbit_r74_c58 bl_58 br_58 wl_74 vdd gnd cell_6t
Xbit_r75_c58 bl_58 br_58 wl_75 vdd gnd cell_6t
Xbit_r76_c58 bl_58 br_58 wl_76 vdd gnd cell_6t
Xbit_r77_c58 bl_58 br_58 wl_77 vdd gnd cell_6t
Xbit_r78_c58 bl_58 br_58 wl_78 vdd gnd cell_6t
Xbit_r79_c58 bl_58 br_58 wl_79 vdd gnd cell_6t
Xbit_r80_c58 bl_58 br_58 wl_80 vdd gnd cell_6t
Xbit_r81_c58 bl_58 br_58 wl_81 vdd gnd cell_6t
Xbit_r82_c58 bl_58 br_58 wl_82 vdd gnd cell_6t
Xbit_r83_c58 bl_58 br_58 wl_83 vdd gnd cell_6t
Xbit_r84_c58 bl_58 br_58 wl_84 vdd gnd cell_6t
Xbit_r85_c58 bl_58 br_58 wl_85 vdd gnd cell_6t
Xbit_r86_c58 bl_58 br_58 wl_86 vdd gnd cell_6t
Xbit_r87_c58 bl_58 br_58 wl_87 vdd gnd cell_6t
Xbit_r88_c58 bl_58 br_58 wl_88 vdd gnd cell_6t
Xbit_r89_c58 bl_58 br_58 wl_89 vdd gnd cell_6t
Xbit_r90_c58 bl_58 br_58 wl_90 vdd gnd cell_6t
Xbit_r91_c58 bl_58 br_58 wl_91 vdd gnd cell_6t
Xbit_r92_c58 bl_58 br_58 wl_92 vdd gnd cell_6t
Xbit_r93_c58 bl_58 br_58 wl_93 vdd gnd cell_6t
Xbit_r94_c58 bl_58 br_58 wl_94 vdd gnd cell_6t
Xbit_r95_c58 bl_58 br_58 wl_95 vdd gnd cell_6t
Xbit_r96_c58 bl_58 br_58 wl_96 vdd gnd cell_6t
Xbit_r97_c58 bl_58 br_58 wl_97 vdd gnd cell_6t
Xbit_r98_c58 bl_58 br_58 wl_98 vdd gnd cell_6t
Xbit_r99_c58 bl_58 br_58 wl_99 vdd gnd cell_6t
Xbit_r100_c58 bl_58 br_58 wl_100 vdd gnd cell_6t
Xbit_r101_c58 bl_58 br_58 wl_101 vdd gnd cell_6t
Xbit_r102_c58 bl_58 br_58 wl_102 vdd gnd cell_6t
Xbit_r103_c58 bl_58 br_58 wl_103 vdd gnd cell_6t
Xbit_r104_c58 bl_58 br_58 wl_104 vdd gnd cell_6t
Xbit_r105_c58 bl_58 br_58 wl_105 vdd gnd cell_6t
Xbit_r106_c58 bl_58 br_58 wl_106 vdd gnd cell_6t
Xbit_r107_c58 bl_58 br_58 wl_107 vdd gnd cell_6t
Xbit_r108_c58 bl_58 br_58 wl_108 vdd gnd cell_6t
Xbit_r109_c58 bl_58 br_58 wl_109 vdd gnd cell_6t
Xbit_r110_c58 bl_58 br_58 wl_110 vdd gnd cell_6t
Xbit_r111_c58 bl_58 br_58 wl_111 vdd gnd cell_6t
Xbit_r112_c58 bl_58 br_58 wl_112 vdd gnd cell_6t
Xbit_r113_c58 bl_58 br_58 wl_113 vdd gnd cell_6t
Xbit_r114_c58 bl_58 br_58 wl_114 vdd gnd cell_6t
Xbit_r115_c58 bl_58 br_58 wl_115 vdd gnd cell_6t
Xbit_r116_c58 bl_58 br_58 wl_116 vdd gnd cell_6t
Xbit_r117_c58 bl_58 br_58 wl_117 vdd gnd cell_6t
Xbit_r118_c58 bl_58 br_58 wl_118 vdd gnd cell_6t
Xbit_r119_c58 bl_58 br_58 wl_119 vdd gnd cell_6t
Xbit_r120_c58 bl_58 br_58 wl_120 vdd gnd cell_6t
Xbit_r121_c58 bl_58 br_58 wl_121 vdd gnd cell_6t
Xbit_r122_c58 bl_58 br_58 wl_122 vdd gnd cell_6t
Xbit_r123_c58 bl_58 br_58 wl_123 vdd gnd cell_6t
Xbit_r124_c58 bl_58 br_58 wl_124 vdd gnd cell_6t
Xbit_r125_c58 bl_58 br_58 wl_125 vdd gnd cell_6t
Xbit_r126_c58 bl_58 br_58 wl_126 vdd gnd cell_6t
Xbit_r127_c58 bl_58 br_58 wl_127 vdd gnd cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd cell_6t
Xbit_r1_c59 bl_59 br_59 wl_1 vdd gnd cell_6t
Xbit_r2_c59 bl_59 br_59 wl_2 vdd gnd cell_6t
Xbit_r3_c59 bl_59 br_59 wl_3 vdd gnd cell_6t
Xbit_r4_c59 bl_59 br_59 wl_4 vdd gnd cell_6t
Xbit_r5_c59 bl_59 br_59 wl_5 vdd gnd cell_6t
Xbit_r6_c59 bl_59 br_59 wl_6 vdd gnd cell_6t
Xbit_r7_c59 bl_59 br_59 wl_7 vdd gnd cell_6t
Xbit_r8_c59 bl_59 br_59 wl_8 vdd gnd cell_6t
Xbit_r9_c59 bl_59 br_59 wl_9 vdd gnd cell_6t
Xbit_r10_c59 bl_59 br_59 wl_10 vdd gnd cell_6t
Xbit_r11_c59 bl_59 br_59 wl_11 vdd gnd cell_6t
Xbit_r12_c59 bl_59 br_59 wl_12 vdd gnd cell_6t
Xbit_r13_c59 bl_59 br_59 wl_13 vdd gnd cell_6t
Xbit_r14_c59 bl_59 br_59 wl_14 vdd gnd cell_6t
Xbit_r15_c59 bl_59 br_59 wl_15 vdd gnd cell_6t
Xbit_r16_c59 bl_59 br_59 wl_16 vdd gnd cell_6t
Xbit_r17_c59 bl_59 br_59 wl_17 vdd gnd cell_6t
Xbit_r18_c59 bl_59 br_59 wl_18 vdd gnd cell_6t
Xbit_r19_c59 bl_59 br_59 wl_19 vdd gnd cell_6t
Xbit_r20_c59 bl_59 br_59 wl_20 vdd gnd cell_6t
Xbit_r21_c59 bl_59 br_59 wl_21 vdd gnd cell_6t
Xbit_r22_c59 bl_59 br_59 wl_22 vdd gnd cell_6t
Xbit_r23_c59 bl_59 br_59 wl_23 vdd gnd cell_6t
Xbit_r24_c59 bl_59 br_59 wl_24 vdd gnd cell_6t
Xbit_r25_c59 bl_59 br_59 wl_25 vdd gnd cell_6t
Xbit_r26_c59 bl_59 br_59 wl_26 vdd gnd cell_6t
Xbit_r27_c59 bl_59 br_59 wl_27 vdd gnd cell_6t
Xbit_r28_c59 bl_59 br_59 wl_28 vdd gnd cell_6t
Xbit_r29_c59 bl_59 br_59 wl_29 vdd gnd cell_6t
Xbit_r30_c59 bl_59 br_59 wl_30 vdd gnd cell_6t
Xbit_r31_c59 bl_59 br_59 wl_31 vdd gnd cell_6t
Xbit_r32_c59 bl_59 br_59 wl_32 vdd gnd cell_6t
Xbit_r33_c59 bl_59 br_59 wl_33 vdd gnd cell_6t
Xbit_r34_c59 bl_59 br_59 wl_34 vdd gnd cell_6t
Xbit_r35_c59 bl_59 br_59 wl_35 vdd gnd cell_6t
Xbit_r36_c59 bl_59 br_59 wl_36 vdd gnd cell_6t
Xbit_r37_c59 bl_59 br_59 wl_37 vdd gnd cell_6t
Xbit_r38_c59 bl_59 br_59 wl_38 vdd gnd cell_6t
Xbit_r39_c59 bl_59 br_59 wl_39 vdd gnd cell_6t
Xbit_r40_c59 bl_59 br_59 wl_40 vdd gnd cell_6t
Xbit_r41_c59 bl_59 br_59 wl_41 vdd gnd cell_6t
Xbit_r42_c59 bl_59 br_59 wl_42 vdd gnd cell_6t
Xbit_r43_c59 bl_59 br_59 wl_43 vdd gnd cell_6t
Xbit_r44_c59 bl_59 br_59 wl_44 vdd gnd cell_6t
Xbit_r45_c59 bl_59 br_59 wl_45 vdd gnd cell_6t
Xbit_r46_c59 bl_59 br_59 wl_46 vdd gnd cell_6t
Xbit_r47_c59 bl_59 br_59 wl_47 vdd gnd cell_6t
Xbit_r48_c59 bl_59 br_59 wl_48 vdd gnd cell_6t
Xbit_r49_c59 bl_59 br_59 wl_49 vdd gnd cell_6t
Xbit_r50_c59 bl_59 br_59 wl_50 vdd gnd cell_6t
Xbit_r51_c59 bl_59 br_59 wl_51 vdd gnd cell_6t
Xbit_r52_c59 bl_59 br_59 wl_52 vdd gnd cell_6t
Xbit_r53_c59 bl_59 br_59 wl_53 vdd gnd cell_6t
Xbit_r54_c59 bl_59 br_59 wl_54 vdd gnd cell_6t
Xbit_r55_c59 bl_59 br_59 wl_55 vdd gnd cell_6t
Xbit_r56_c59 bl_59 br_59 wl_56 vdd gnd cell_6t
Xbit_r57_c59 bl_59 br_59 wl_57 vdd gnd cell_6t
Xbit_r58_c59 bl_59 br_59 wl_58 vdd gnd cell_6t
Xbit_r59_c59 bl_59 br_59 wl_59 vdd gnd cell_6t
Xbit_r60_c59 bl_59 br_59 wl_60 vdd gnd cell_6t
Xbit_r61_c59 bl_59 br_59 wl_61 vdd gnd cell_6t
Xbit_r62_c59 bl_59 br_59 wl_62 vdd gnd cell_6t
Xbit_r63_c59 bl_59 br_59 wl_63 vdd gnd cell_6t
Xbit_r64_c59 bl_59 br_59 wl_64 vdd gnd cell_6t
Xbit_r65_c59 bl_59 br_59 wl_65 vdd gnd cell_6t
Xbit_r66_c59 bl_59 br_59 wl_66 vdd gnd cell_6t
Xbit_r67_c59 bl_59 br_59 wl_67 vdd gnd cell_6t
Xbit_r68_c59 bl_59 br_59 wl_68 vdd gnd cell_6t
Xbit_r69_c59 bl_59 br_59 wl_69 vdd gnd cell_6t
Xbit_r70_c59 bl_59 br_59 wl_70 vdd gnd cell_6t
Xbit_r71_c59 bl_59 br_59 wl_71 vdd gnd cell_6t
Xbit_r72_c59 bl_59 br_59 wl_72 vdd gnd cell_6t
Xbit_r73_c59 bl_59 br_59 wl_73 vdd gnd cell_6t
Xbit_r74_c59 bl_59 br_59 wl_74 vdd gnd cell_6t
Xbit_r75_c59 bl_59 br_59 wl_75 vdd gnd cell_6t
Xbit_r76_c59 bl_59 br_59 wl_76 vdd gnd cell_6t
Xbit_r77_c59 bl_59 br_59 wl_77 vdd gnd cell_6t
Xbit_r78_c59 bl_59 br_59 wl_78 vdd gnd cell_6t
Xbit_r79_c59 bl_59 br_59 wl_79 vdd gnd cell_6t
Xbit_r80_c59 bl_59 br_59 wl_80 vdd gnd cell_6t
Xbit_r81_c59 bl_59 br_59 wl_81 vdd gnd cell_6t
Xbit_r82_c59 bl_59 br_59 wl_82 vdd gnd cell_6t
Xbit_r83_c59 bl_59 br_59 wl_83 vdd gnd cell_6t
Xbit_r84_c59 bl_59 br_59 wl_84 vdd gnd cell_6t
Xbit_r85_c59 bl_59 br_59 wl_85 vdd gnd cell_6t
Xbit_r86_c59 bl_59 br_59 wl_86 vdd gnd cell_6t
Xbit_r87_c59 bl_59 br_59 wl_87 vdd gnd cell_6t
Xbit_r88_c59 bl_59 br_59 wl_88 vdd gnd cell_6t
Xbit_r89_c59 bl_59 br_59 wl_89 vdd gnd cell_6t
Xbit_r90_c59 bl_59 br_59 wl_90 vdd gnd cell_6t
Xbit_r91_c59 bl_59 br_59 wl_91 vdd gnd cell_6t
Xbit_r92_c59 bl_59 br_59 wl_92 vdd gnd cell_6t
Xbit_r93_c59 bl_59 br_59 wl_93 vdd gnd cell_6t
Xbit_r94_c59 bl_59 br_59 wl_94 vdd gnd cell_6t
Xbit_r95_c59 bl_59 br_59 wl_95 vdd gnd cell_6t
Xbit_r96_c59 bl_59 br_59 wl_96 vdd gnd cell_6t
Xbit_r97_c59 bl_59 br_59 wl_97 vdd gnd cell_6t
Xbit_r98_c59 bl_59 br_59 wl_98 vdd gnd cell_6t
Xbit_r99_c59 bl_59 br_59 wl_99 vdd gnd cell_6t
Xbit_r100_c59 bl_59 br_59 wl_100 vdd gnd cell_6t
Xbit_r101_c59 bl_59 br_59 wl_101 vdd gnd cell_6t
Xbit_r102_c59 bl_59 br_59 wl_102 vdd gnd cell_6t
Xbit_r103_c59 bl_59 br_59 wl_103 vdd gnd cell_6t
Xbit_r104_c59 bl_59 br_59 wl_104 vdd gnd cell_6t
Xbit_r105_c59 bl_59 br_59 wl_105 vdd gnd cell_6t
Xbit_r106_c59 bl_59 br_59 wl_106 vdd gnd cell_6t
Xbit_r107_c59 bl_59 br_59 wl_107 vdd gnd cell_6t
Xbit_r108_c59 bl_59 br_59 wl_108 vdd gnd cell_6t
Xbit_r109_c59 bl_59 br_59 wl_109 vdd gnd cell_6t
Xbit_r110_c59 bl_59 br_59 wl_110 vdd gnd cell_6t
Xbit_r111_c59 bl_59 br_59 wl_111 vdd gnd cell_6t
Xbit_r112_c59 bl_59 br_59 wl_112 vdd gnd cell_6t
Xbit_r113_c59 bl_59 br_59 wl_113 vdd gnd cell_6t
Xbit_r114_c59 bl_59 br_59 wl_114 vdd gnd cell_6t
Xbit_r115_c59 bl_59 br_59 wl_115 vdd gnd cell_6t
Xbit_r116_c59 bl_59 br_59 wl_116 vdd gnd cell_6t
Xbit_r117_c59 bl_59 br_59 wl_117 vdd gnd cell_6t
Xbit_r118_c59 bl_59 br_59 wl_118 vdd gnd cell_6t
Xbit_r119_c59 bl_59 br_59 wl_119 vdd gnd cell_6t
Xbit_r120_c59 bl_59 br_59 wl_120 vdd gnd cell_6t
Xbit_r121_c59 bl_59 br_59 wl_121 vdd gnd cell_6t
Xbit_r122_c59 bl_59 br_59 wl_122 vdd gnd cell_6t
Xbit_r123_c59 bl_59 br_59 wl_123 vdd gnd cell_6t
Xbit_r124_c59 bl_59 br_59 wl_124 vdd gnd cell_6t
Xbit_r125_c59 bl_59 br_59 wl_125 vdd gnd cell_6t
Xbit_r126_c59 bl_59 br_59 wl_126 vdd gnd cell_6t
Xbit_r127_c59 bl_59 br_59 wl_127 vdd gnd cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd cell_6t
Xbit_r1_c60 bl_60 br_60 wl_1 vdd gnd cell_6t
Xbit_r2_c60 bl_60 br_60 wl_2 vdd gnd cell_6t
Xbit_r3_c60 bl_60 br_60 wl_3 vdd gnd cell_6t
Xbit_r4_c60 bl_60 br_60 wl_4 vdd gnd cell_6t
Xbit_r5_c60 bl_60 br_60 wl_5 vdd gnd cell_6t
Xbit_r6_c60 bl_60 br_60 wl_6 vdd gnd cell_6t
Xbit_r7_c60 bl_60 br_60 wl_7 vdd gnd cell_6t
Xbit_r8_c60 bl_60 br_60 wl_8 vdd gnd cell_6t
Xbit_r9_c60 bl_60 br_60 wl_9 vdd gnd cell_6t
Xbit_r10_c60 bl_60 br_60 wl_10 vdd gnd cell_6t
Xbit_r11_c60 bl_60 br_60 wl_11 vdd gnd cell_6t
Xbit_r12_c60 bl_60 br_60 wl_12 vdd gnd cell_6t
Xbit_r13_c60 bl_60 br_60 wl_13 vdd gnd cell_6t
Xbit_r14_c60 bl_60 br_60 wl_14 vdd gnd cell_6t
Xbit_r15_c60 bl_60 br_60 wl_15 vdd gnd cell_6t
Xbit_r16_c60 bl_60 br_60 wl_16 vdd gnd cell_6t
Xbit_r17_c60 bl_60 br_60 wl_17 vdd gnd cell_6t
Xbit_r18_c60 bl_60 br_60 wl_18 vdd gnd cell_6t
Xbit_r19_c60 bl_60 br_60 wl_19 vdd gnd cell_6t
Xbit_r20_c60 bl_60 br_60 wl_20 vdd gnd cell_6t
Xbit_r21_c60 bl_60 br_60 wl_21 vdd gnd cell_6t
Xbit_r22_c60 bl_60 br_60 wl_22 vdd gnd cell_6t
Xbit_r23_c60 bl_60 br_60 wl_23 vdd gnd cell_6t
Xbit_r24_c60 bl_60 br_60 wl_24 vdd gnd cell_6t
Xbit_r25_c60 bl_60 br_60 wl_25 vdd gnd cell_6t
Xbit_r26_c60 bl_60 br_60 wl_26 vdd gnd cell_6t
Xbit_r27_c60 bl_60 br_60 wl_27 vdd gnd cell_6t
Xbit_r28_c60 bl_60 br_60 wl_28 vdd gnd cell_6t
Xbit_r29_c60 bl_60 br_60 wl_29 vdd gnd cell_6t
Xbit_r30_c60 bl_60 br_60 wl_30 vdd gnd cell_6t
Xbit_r31_c60 bl_60 br_60 wl_31 vdd gnd cell_6t
Xbit_r32_c60 bl_60 br_60 wl_32 vdd gnd cell_6t
Xbit_r33_c60 bl_60 br_60 wl_33 vdd gnd cell_6t
Xbit_r34_c60 bl_60 br_60 wl_34 vdd gnd cell_6t
Xbit_r35_c60 bl_60 br_60 wl_35 vdd gnd cell_6t
Xbit_r36_c60 bl_60 br_60 wl_36 vdd gnd cell_6t
Xbit_r37_c60 bl_60 br_60 wl_37 vdd gnd cell_6t
Xbit_r38_c60 bl_60 br_60 wl_38 vdd gnd cell_6t
Xbit_r39_c60 bl_60 br_60 wl_39 vdd gnd cell_6t
Xbit_r40_c60 bl_60 br_60 wl_40 vdd gnd cell_6t
Xbit_r41_c60 bl_60 br_60 wl_41 vdd gnd cell_6t
Xbit_r42_c60 bl_60 br_60 wl_42 vdd gnd cell_6t
Xbit_r43_c60 bl_60 br_60 wl_43 vdd gnd cell_6t
Xbit_r44_c60 bl_60 br_60 wl_44 vdd gnd cell_6t
Xbit_r45_c60 bl_60 br_60 wl_45 vdd gnd cell_6t
Xbit_r46_c60 bl_60 br_60 wl_46 vdd gnd cell_6t
Xbit_r47_c60 bl_60 br_60 wl_47 vdd gnd cell_6t
Xbit_r48_c60 bl_60 br_60 wl_48 vdd gnd cell_6t
Xbit_r49_c60 bl_60 br_60 wl_49 vdd gnd cell_6t
Xbit_r50_c60 bl_60 br_60 wl_50 vdd gnd cell_6t
Xbit_r51_c60 bl_60 br_60 wl_51 vdd gnd cell_6t
Xbit_r52_c60 bl_60 br_60 wl_52 vdd gnd cell_6t
Xbit_r53_c60 bl_60 br_60 wl_53 vdd gnd cell_6t
Xbit_r54_c60 bl_60 br_60 wl_54 vdd gnd cell_6t
Xbit_r55_c60 bl_60 br_60 wl_55 vdd gnd cell_6t
Xbit_r56_c60 bl_60 br_60 wl_56 vdd gnd cell_6t
Xbit_r57_c60 bl_60 br_60 wl_57 vdd gnd cell_6t
Xbit_r58_c60 bl_60 br_60 wl_58 vdd gnd cell_6t
Xbit_r59_c60 bl_60 br_60 wl_59 vdd gnd cell_6t
Xbit_r60_c60 bl_60 br_60 wl_60 vdd gnd cell_6t
Xbit_r61_c60 bl_60 br_60 wl_61 vdd gnd cell_6t
Xbit_r62_c60 bl_60 br_60 wl_62 vdd gnd cell_6t
Xbit_r63_c60 bl_60 br_60 wl_63 vdd gnd cell_6t
Xbit_r64_c60 bl_60 br_60 wl_64 vdd gnd cell_6t
Xbit_r65_c60 bl_60 br_60 wl_65 vdd gnd cell_6t
Xbit_r66_c60 bl_60 br_60 wl_66 vdd gnd cell_6t
Xbit_r67_c60 bl_60 br_60 wl_67 vdd gnd cell_6t
Xbit_r68_c60 bl_60 br_60 wl_68 vdd gnd cell_6t
Xbit_r69_c60 bl_60 br_60 wl_69 vdd gnd cell_6t
Xbit_r70_c60 bl_60 br_60 wl_70 vdd gnd cell_6t
Xbit_r71_c60 bl_60 br_60 wl_71 vdd gnd cell_6t
Xbit_r72_c60 bl_60 br_60 wl_72 vdd gnd cell_6t
Xbit_r73_c60 bl_60 br_60 wl_73 vdd gnd cell_6t
Xbit_r74_c60 bl_60 br_60 wl_74 vdd gnd cell_6t
Xbit_r75_c60 bl_60 br_60 wl_75 vdd gnd cell_6t
Xbit_r76_c60 bl_60 br_60 wl_76 vdd gnd cell_6t
Xbit_r77_c60 bl_60 br_60 wl_77 vdd gnd cell_6t
Xbit_r78_c60 bl_60 br_60 wl_78 vdd gnd cell_6t
Xbit_r79_c60 bl_60 br_60 wl_79 vdd gnd cell_6t
Xbit_r80_c60 bl_60 br_60 wl_80 vdd gnd cell_6t
Xbit_r81_c60 bl_60 br_60 wl_81 vdd gnd cell_6t
Xbit_r82_c60 bl_60 br_60 wl_82 vdd gnd cell_6t
Xbit_r83_c60 bl_60 br_60 wl_83 vdd gnd cell_6t
Xbit_r84_c60 bl_60 br_60 wl_84 vdd gnd cell_6t
Xbit_r85_c60 bl_60 br_60 wl_85 vdd gnd cell_6t
Xbit_r86_c60 bl_60 br_60 wl_86 vdd gnd cell_6t
Xbit_r87_c60 bl_60 br_60 wl_87 vdd gnd cell_6t
Xbit_r88_c60 bl_60 br_60 wl_88 vdd gnd cell_6t
Xbit_r89_c60 bl_60 br_60 wl_89 vdd gnd cell_6t
Xbit_r90_c60 bl_60 br_60 wl_90 vdd gnd cell_6t
Xbit_r91_c60 bl_60 br_60 wl_91 vdd gnd cell_6t
Xbit_r92_c60 bl_60 br_60 wl_92 vdd gnd cell_6t
Xbit_r93_c60 bl_60 br_60 wl_93 vdd gnd cell_6t
Xbit_r94_c60 bl_60 br_60 wl_94 vdd gnd cell_6t
Xbit_r95_c60 bl_60 br_60 wl_95 vdd gnd cell_6t
Xbit_r96_c60 bl_60 br_60 wl_96 vdd gnd cell_6t
Xbit_r97_c60 bl_60 br_60 wl_97 vdd gnd cell_6t
Xbit_r98_c60 bl_60 br_60 wl_98 vdd gnd cell_6t
Xbit_r99_c60 bl_60 br_60 wl_99 vdd gnd cell_6t
Xbit_r100_c60 bl_60 br_60 wl_100 vdd gnd cell_6t
Xbit_r101_c60 bl_60 br_60 wl_101 vdd gnd cell_6t
Xbit_r102_c60 bl_60 br_60 wl_102 vdd gnd cell_6t
Xbit_r103_c60 bl_60 br_60 wl_103 vdd gnd cell_6t
Xbit_r104_c60 bl_60 br_60 wl_104 vdd gnd cell_6t
Xbit_r105_c60 bl_60 br_60 wl_105 vdd gnd cell_6t
Xbit_r106_c60 bl_60 br_60 wl_106 vdd gnd cell_6t
Xbit_r107_c60 bl_60 br_60 wl_107 vdd gnd cell_6t
Xbit_r108_c60 bl_60 br_60 wl_108 vdd gnd cell_6t
Xbit_r109_c60 bl_60 br_60 wl_109 vdd gnd cell_6t
Xbit_r110_c60 bl_60 br_60 wl_110 vdd gnd cell_6t
Xbit_r111_c60 bl_60 br_60 wl_111 vdd gnd cell_6t
Xbit_r112_c60 bl_60 br_60 wl_112 vdd gnd cell_6t
Xbit_r113_c60 bl_60 br_60 wl_113 vdd gnd cell_6t
Xbit_r114_c60 bl_60 br_60 wl_114 vdd gnd cell_6t
Xbit_r115_c60 bl_60 br_60 wl_115 vdd gnd cell_6t
Xbit_r116_c60 bl_60 br_60 wl_116 vdd gnd cell_6t
Xbit_r117_c60 bl_60 br_60 wl_117 vdd gnd cell_6t
Xbit_r118_c60 bl_60 br_60 wl_118 vdd gnd cell_6t
Xbit_r119_c60 bl_60 br_60 wl_119 vdd gnd cell_6t
Xbit_r120_c60 bl_60 br_60 wl_120 vdd gnd cell_6t
Xbit_r121_c60 bl_60 br_60 wl_121 vdd gnd cell_6t
Xbit_r122_c60 bl_60 br_60 wl_122 vdd gnd cell_6t
Xbit_r123_c60 bl_60 br_60 wl_123 vdd gnd cell_6t
Xbit_r124_c60 bl_60 br_60 wl_124 vdd gnd cell_6t
Xbit_r125_c60 bl_60 br_60 wl_125 vdd gnd cell_6t
Xbit_r126_c60 bl_60 br_60 wl_126 vdd gnd cell_6t
Xbit_r127_c60 bl_60 br_60 wl_127 vdd gnd cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd cell_6t
Xbit_r1_c61 bl_61 br_61 wl_1 vdd gnd cell_6t
Xbit_r2_c61 bl_61 br_61 wl_2 vdd gnd cell_6t
Xbit_r3_c61 bl_61 br_61 wl_3 vdd gnd cell_6t
Xbit_r4_c61 bl_61 br_61 wl_4 vdd gnd cell_6t
Xbit_r5_c61 bl_61 br_61 wl_5 vdd gnd cell_6t
Xbit_r6_c61 bl_61 br_61 wl_6 vdd gnd cell_6t
Xbit_r7_c61 bl_61 br_61 wl_7 vdd gnd cell_6t
Xbit_r8_c61 bl_61 br_61 wl_8 vdd gnd cell_6t
Xbit_r9_c61 bl_61 br_61 wl_9 vdd gnd cell_6t
Xbit_r10_c61 bl_61 br_61 wl_10 vdd gnd cell_6t
Xbit_r11_c61 bl_61 br_61 wl_11 vdd gnd cell_6t
Xbit_r12_c61 bl_61 br_61 wl_12 vdd gnd cell_6t
Xbit_r13_c61 bl_61 br_61 wl_13 vdd gnd cell_6t
Xbit_r14_c61 bl_61 br_61 wl_14 vdd gnd cell_6t
Xbit_r15_c61 bl_61 br_61 wl_15 vdd gnd cell_6t
Xbit_r16_c61 bl_61 br_61 wl_16 vdd gnd cell_6t
Xbit_r17_c61 bl_61 br_61 wl_17 vdd gnd cell_6t
Xbit_r18_c61 bl_61 br_61 wl_18 vdd gnd cell_6t
Xbit_r19_c61 bl_61 br_61 wl_19 vdd gnd cell_6t
Xbit_r20_c61 bl_61 br_61 wl_20 vdd gnd cell_6t
Xbit_r21_c61 bl_61 br_61 wl_21 vdd gnd cell_6t
Xbit_r22_c61 bl_61 br_61 wl_22 vdd gnd cell_6t
Xbit_r23_c61 bl_61 br_61 wl_23 vdd gnd cell_6t
Xbit_r24_c61 bl_61 br_61 wl_24 vdd gnd cell_6t
Xbit_r25_c61 bl_61 br_61 wl_25 vdd gnd cell_6t
Xbit_r26_c61 bl_61 br_61 wl_26 vdd gnd cell_6t
Xbit_r27_c61 bl_61 br_61 wl_27 vdd gnd cell_6t
Xbit_r28_c61 bl_61 br_61 wl_28 vdd gnd cell_6t
Xbit_r29_c61 bl_61 br_61 wl_29 vdd gnd cell_6t
Xbit_r30_c61 bl_61 br_61 wl_30 vdd gnd cell_6t
Xbit_r31_c61 bl_61 br_61 wl_31 vdd gnd cell_6t
Xbit_r32_c61 bl_61 br_61 wl_32 vdd gnd cell_6t
Xbit_r33_c61 bl_61 br_61 wl_33 vdd gnd cell_6t
Xbit_r34_c61 bl_61 br_61 wl_34 vdd gnd cell_6t
Xbit_r35_c61 bl_61 br_61 wl_35 vdd gnd cell_6t
Xbit_r36_c61 bl_61 br_61 wl_36 vdd gnd cell_6t
Xbit_r37_c61 bl_61 br_61 wl_37 vdd gnd cell_6t
Xbit_r38_c61 bl_61 br_61 wl_38 vdd gnd cell_6t
Xbit_r39_c61 bl_61 br_61 wl_39 vdd gnd cell_6t
Xbit_r40_c61 bl_61 br_61 wl_40 vdd gnd cell_6t
Xbit_r41_c61 bl_61 br_61 wl_41 vdd gnd cell_6t
Xbit_r42_c61 bl_61 br_61 wl_42 vdd gnd cell_6t
Xbit_r43_c61 bl_61 br_61 wl_43 vdd gnd cell_6t
Xbit_r44_c61 bl_61 br_61 wl_44 vdd gnd cell_6t
Xbit_r45_c61 bl_61 br_61 wl_45 vdd gnd cell_6t
Xbit_r46_c61 bl_61 br_61 wl_46 vdd gnd cell_6t
Xbit_r47_c61 bl_61 br_61 wl_47 vdd gnd cell_6t
Xbit_r48_c61 bl_61 br_61 wl_48 vdd gnd cell_6t
Xbit_r49_c61 bl_61 br_61 wl_49 vdd gnd cell_6t
Xbit_r50_c61 bl_61 br_61 wl_50 vdd gnd cell_6t
Xbit_r51_c61 bl_61 br_61 wl_51 vdd gnd cell_6t
Xbit_r52_c61 bl_61 br_61 wl_52 vdd gnd cell_6t
Xbit_r53_c61 bl_61 br_61 wl_53 vdd gnd cell_6t
Xbit_r54_c61 bl_61 br_61 wl_54 vdd gnd cell_6t
Xbit_r55_c61 bl_61 br_61 wl_55 vdd gnd cell_6t
Xbit_r56_c61 bl_61 br_61 wl_56 vdd gnd cell_6t
Xbit_r57_c61 bl_61 br_61 wl_57 vdd gnd cell_6t
Xbit_r58_c61 bl_61 br_61 wl_58 vdd gnd cell_6t
Xbit_r59_c61 bl_61 br_61 wl_59 vdd gnd cell_6t
Xbit_r60_c61 bl_61 br_61 wl_60 vdd gnd cell_6t
Xbit_r61_c61 bl_61 br_61 wl_61 vdd gnd cell_6t
Xbit_r62_c61 bl_61 br_61 wl_62 vdd gnd cell_6t
Xbit_r63_c61 bl_61 br_61 wl_63 vdd gnd cell_6t
Xbit_r64_c61 bl_61 br_61 wl_64 vdd gnd cell_6t
Xbit_r65_c61 bl_61 br_61 wl_65 vdd gnd cell_6t
Xbit_r66_c61 bl_61 br_61 wl_66 vdd gnd cell_6t
Xbit_r67_c61 bl_61 br_61 wl_67 vdd gnd cell_6t
Xbit_r68_c61 bl_61 br_61 wl_68 vdd gnd cell_6t
Xbit_r69_c61 bl_61 br_61 wl_69 vdd gnd cell_6t
Xbit_r70_c61 bl_61 br_61 wl_70 vdd gnd cell_6t
Xbit_r71_c61 bl_61 br_61 wl_71 vdd gnd cell_6t
Xbit_r72_c61 bl_61 br_61 wl_72 vdd gnd cell_6t
Xbit_r73_c61 bl_61 br_61 wl_73 vdd gnd cell_6t
Xbit_r74_c61 bl_61 br_61 wl_74 vdd gnd cell_6t
Xbit_r75_c61 bl_61 br_61 wl_75 vdd gnd cell_6t
Xbit_r76_c61 bl_61 br_61 wl_76 vdd gnd cell_6t
Xbit_r77_c61 bl_61 br_61 wl_77 vdd gnd cell_6t
Xbit_r78_c61 bl_61 br_61 wl_78 vdd gnd cell_6t
Xbit_r79_c61 bl_61 br_61 wl_79 vdd gnd cell_6t
Xbit_r80_c61 bl_61 br_61 wl_80 vdd gnd cell_6t
Xbit_r81_c61 bl_61 br_61 wl_81 vdd gnd cell_6t
Xbit_r82_c61 bl_61 br_61 wl_82 vdd gnd cell_6t
Xbit_r83_c61 bl_61 br_61 wl_83 vdd gnd cell_6t
Xbit_r84_c61 bl_61 br_61 wl_84 vdd gnd cell_6t
Xbit_r85_c61 bl_61 br_61 wl_85 vdd gnd cell_6t
Xbit_r86_c61 bl_61 br_61 wl_86 vdd gnd cell_6t
Xbit_r87_c61 bl_61 br_61 wl_87 vdd gnd cell_6t
Xbit_r88_c61 bl_61 br_61 wl_88 vdd gnd cell_6t
Xbit_r89_c61 bl_61 br_61 wl_89 vdd gnd cell_6t
Xbit_r90_c61 bl_61 br_61 wl_90 vdd gnd cell_6t
Xbit_r91_c61 bl_61 br_61 wl_91 vdd gnd cell_6t
Xbit_r92_c61 bl_61 br_61 wl_92 vdd gnd cell_6t
Xbit_r93_c61 bl_61 br_61 wl_93 vdd gnd cell_6t
Xbit_r94_c61 bl_61 br_61 wl_94 vdd gnd cell_6t
Xbit_r95_c61 bl_61 br_61 wl_95 vdd gnd cell_6t
Xbit_r96_c61 bl_61 br_61 wl_96 vdd gnd cell_6t
Xbit_r97_c61 bl_61 br_61 wl_97 vdd gnd cell_6t
Xbit_r98_c61 bl_61 br_61 wl_98 vdd gnd cell_6t
Xbit_r99_c61 bl_61 br_61 wl_99 vdd gnd cell_6t
Xbit_r100_c61 bl_61 br_61 wl_100 vdd gnd cell_6t
Xbit_r101_c61 bl_61 br_61 wl_101 vdd gnd cell_6t
Xbit_r102_c61 bl_61 br_61 wl_102 vdd gnd cell_6t
Xbit_r103_c61 bl_61 br_61 wl_103 vdd gnd cell_6t
Xbit_r104_c61 bl_61 br_61 wl_104 vdd gnd cell_6t
Xbit_r105_c61 bl_61 br_61 wl_105 vdd gnd cell_6t
Xbit_r106_c61 bl_61 br_61 wl_106 vdd gnd cell_6t
Xbit_r107_c61 bl_61 br_61 wl_107 vdd gnd cell_6t
Xbit_r108_c61 bl_61 br_61 wl_108 vdd gnd cell_6t
Xbit_r109_c61 bl_61 br_61 wl_109 vdd gnd cell_6t
Xbit_r110_c61 bl_61 br_61 wl_110 vdd gnd cell_6t
Xbit_r111_c61 bl_61 br_61 wl_111 vdd gnd cell_6t
Xbit_r112_c61 bl_61 br_61 wl_112 vdd gnd cell_6t
Xbit_r113_c61 bl_61 br_61 wl_113 vdd gnd cell_6t
Xbit_r114_c61 bl_61 br_61 wl_114 vdd gnd cell_6t
Xbit_r115_c61 bl_61 br_61 wl_115 vdd gnd cell_6t
Xbit_r116_c61 bl_61 br_61 wl_116 vdd gnd cell_6t
Xbit_r117_c61 bl_61 br_61 wl_117 vdd gnd cell_6t
Xbit_r118_c61 bl_61 br_61 wl_118 vdd gnd cell_6t
Xbit_r119_c61 bl_61 br_61 wl_119 vdd gnd cell_6t
Xbit_r120_c61 bl_61 br_61 wl_120 vdd gnd cell_6t
Xbit_r121_c61 bl_61 br_61 wl_121 vdd gnd cell_6t
Xbit_r122_c61 bl_61 br_61 wl_122 vdd gnd cell_6t
Xbit_r123_c61 bl_61 br_61 wl_123 vdd gnd cell_6t
Xbit_r124_c61 bl_61 br_61 wl_124 vdd gnd cell_6t
Xbit_r125_c61 bl_61 br_61 wl_125 vdd gnd cell_6t
Xbit_r126_c61 bl_61 br_61 wl_126 vdd gnd cell_6t
Xbit_r127_c61 bl_61 br_61 wl_127 vdd gnd cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd cell_6t
Xbit_r1_c62 bl_62 br_62 wl_1 vdd gnd cell_6t
Xbit_r2_c62 bl_62 br_62 wl_2 vdd gnd cell_6t
Xbit_r3_c62 bl_62 br_62 wl_3 vdd gnd cell_6t
Xbit_r4_c62 bl_62 br_62 wl_4 vdd gnd cell_6t
Xbit_r5_c62 bl_62 br_62 wl_5 vdd gnd cell_6t
Xbit_r6_c62 bl_62 br_62 wl_6 vdd gnd cell_6t
Xbit_r7_c62 bl_62 br_62 wl_7 vdd gnd cell_6t
Xbit_r8_c62 bl_62 br_62 wl_8 vdd gnd cell_6t
Xbit_r9_c62 bl_62 br_62 wl_9 vdd gnd cell_6t
Xbit_r10_c62 bl_62 br_62 wl_10 vdd gnd cell_6t
Xbit_r11_c62 bl_62 br_62 wl_11 vdd gnd cell_6t
Xbit_r12_c62 bl_62 br_62 wl_12 vdd gnd cell_6t
Xbit_r13_c62 bl_62 br_62 wl_13 vdd gnd cell_6t
Xbit_r14_c62 bl_62 br_62 wl_14 vdd gnd cell_6t
Xbit_r15_c62 bl_62 br_62 wl_15 vdd gnd cell_6t
Xbit_r16_c62 bl_62 br_62 wl_16 vdd gnd cell_6t
Xbit_r17_c62 bl_62 br_62 wl_17 vdd gnd cell_6t
Xbit_r18_c62 bl_62 br_62 wl_18 vdd gnd cell_6t
Xbit_r19_c62 bl_62 br_62 wl_19 vdd gnd cell_6t
Xbit_r20_c62 bl_62 br_62 wl_20 vdd gnd cell_6t
Xbit_r21_c62 bl_62 br_62 wl_21 vdd gnd cell_6t
Xbit_r22_c62 bl_62 br_62 wl_22 vdd gnd cell_6t
Xbit_r23_c62 bl_62 br_62 wl_23 vdd gnd cell_6t
Xbit_r24_c62 bl_62 br_62 wl_24 vdd gnd cell_6t
Xbit_r25_c62 bl_62 br_62 wl_25 vdd gnd cell_6t
Xbit_r26_c62 bl_62 br_62 wl_26 vdd gnd cell_6t
Xbit_r27_c62 bl_62 br_62 wl_27 vdd gnd cell_6t
Xbit_r28_c62 bl_62 br_62 wl_28 vdd gnd cell_6t
Xbit_r29_c62 bl_62 br_62 wl_29 vdd gnd cell_6t
Xbit_r30_c62 bl_62 br_62 wl_30 vdd gnd cell_6t
Xbit_r31_c62 bl_62 br_62 wl_31 vdd gnd cell_6t
Xbit_r32_c62 bl_62 br_62 wl_32 vdd gnd cell_6t
Xbit_r33_c62 bl_62 br_62 wl_33 vdd gnd cell_6t
Xbit_r34_c62 bl_62 br_62 wl_34 vdd gnd cell_6t
Xbit_r35_c62 bl_62 br_62 wl_35 vdd gnd cell_6t
Xbit_r36_c62 bl_62 br_62 wl_36 vdd gnd cell_6t
Xbit_r37_c62 bl_62 br_62 wl_37 vdd gnd cell_6t
Xbit_r38_c62 bl_62 br_62 wl_38 vdd gnd cell_6t
Xbit_r39_c62 bl_62 br_62 wl_39 vdd gnd cell_6t
Xbit_r40_c62 bl_62 br_62 wl_40 vdd gnd cell_6t
Xbit_r41_c62 bl_62 br_62 wl_41 vdd gnd cell_6t
Xbit_r42_c62 bl_62 br_62 wl_42 vdd gnd cell_6t
Xbit_r43_c62 bl_62 br_62 wl_43 vdd gnd cell_6t
Xbit_r44_c62 bl_62 br_62 wl_44 vdd gnd cell_6t
Xbit_r45_c62 bl_62 br_62 wl_45 vdd gnd cell_6t
Xbit_r46_c62 bl_62 br_62 wl_46 vdd gnd cell_6t
Xbit_r47_c62 bl_62 br_62 wl_47 vdd gnd cell_6t
Xbit_r48_c62 bl_62 br_62 wl_48 vdd gnd cell_6t
Xbit_r49_c62 bl_62 br_62 wl_49 vdd gnd cell_6t
Xbit_r50_c62 bl_62 br_62 wl_50 vdd gnd cell_6t
Xbit_r51_c62 bl_62 br_62 wl_51 vdd gnd cell_6t
Xbit_r52_c62 bl_62 br_62 wl_52 vdd gnd cell_6t
Xbit_r53_c62 bl_62 br_62 wl_53 vdd gnd cell_6t
Xbit_r54_c62 bl_62 br_62 wl_54 vdd gnd cell_6t
Xbit_r55_c62 bl_62 br_62 wl_55 vdd gnd cell_6t
Xbit_r56_c62 bl_62 br_62 wl_56 vdd gnd cell_6t
Xbit_r57_c62 bl_62 br_62 wl_57 vdd gnd cell_6t
Xbit_r58_c62 bl_62 br_62 wl_58 vdd gnd cell_6t
Xbit_r59_c62 bl_62 br_62 wl_59 vdd gnd cell_6t
Xbit_r60_c62 bl_62 br_62 wl_60 vdd gnd cell_6t
Xbit_r61_c62 bl_62 br_62 wl_61 vdd gnd cell_6t
Xbit_r62_c62 bl_62 br_62 wl_62 vdd gnd cell_6t
Xbit_r63_c62 bl_62 br_62 wl_63 vdd gnd cell_6t
Xbit_r64_c62 bl_62 br_62 wl_64 vdd gnd cell_6t
Xbit_r65_c62 bl_62 br_62 wl_65 vdd gnd cell_6t
Xbit_r66_c62 bl_62 br_62 wl_66 vdd gnd cell_6t
Xbit_r67_c62 bl_62 br_62 wl_67 vdd gnd cell_6t
Xbit_r68_c62 bl_62 br_62 wl_68 vdd gnd cell_6t
Xbit_r69_c62 bl_62 br_62 wl_69 vdd gnd cell_6t
Xbit_r70_c62 bl_62 br_62 wl_70 vdd gnd cell_6t
Xbit_r71_c62 bl_62 br_62 wl_71 vdd gnd cell_6t
Xbit_r72_c62 bl_62 br_62 wl_72 vdd gnd cell_6t
Xbit_r73_c62 bl_62 br_62 wl_73 vdd gnd cell_6t
Xbit_r74_c62 bl_62 br_62 wl_74 vdd gnd cell_6t
Xbit_r75_c62 bl_62 br_62 wl_75 vdd gnd cell_6t
Xbit_r76_c62 bl_62 br_62 wl_76 vdd gnd cell_6t
Xbit_r77_c62 bl_62 br_62 wl_77 vdd gnd cell_6t
Xbit_r78_c62 bl_62 br_62 wl_78 vdd gnd cell_6t
Xbit_r79_c62 bl_62 br_62 wl_79 vdd gnd cell_6t
Xbit_r80_c62 bl_62 br_62 wl_80 vdd gnd cell_6t
Xbit_r81_c62 bl_62 br_62 wl_81 vdd gnd cell_6t
Xbit_r82_c62 bl_62 br_62 wl_82 vdd gnd cell_6t
Xbit_r83_c62 bl_62 br_62 wl_83 vdd gnd cell_6t
Xbit_r84_c62 bl_62 br_62 wl_84 vdd gnd cell_6t
Xbit_r85_c62 bl_62 br_62 wl_85 vdd gnd cell_6t
Xbit_r86_c62 bl_62 br_62 wl_86 vdd gnd cell_6t
Xbit_r87_c62 bl_62 br_62 wl_87 vdd gnd cell_6t
Xbit_r88_c62 bl_62 br_62 wl_88 vdd gnd cell_6t
Xbit_r89_c62 bl_62 br_62 wl_89 vdd gnd cell_6t
Xbit_r90_c62 bl_62 br_62 wl_90 vdd gnd cell_6t
Xbit_r91_c62 bl_62 br_62 wl_91 vdd gnd cell_6t
Xbit_r92_c62 bl_62 br_62 wl_92 vdd gnd cell_6t
Xbit_r93_c62 bl_62 br_62 wl_93 vdd gnd cell_6t
Xbit_r94_c62 bl_62 br_62 wl_94 vdd gnd cell_6t
Xbit_r95_c62 bl_62 br_62 wl_95 vdd gnd cell_6t
Xbit_r96_c62 bl_62 br_62 wl_96 vdd gnd cell_6t
Xbit_r97_c62 bl_62 br_62 wl_97 vdd gnd cell_6t
Xbit_r98_c62 bl_62 br_62 wl_98 vdd gnd cell_6t
Xbit_r99_c62 bl_62 br_62 wl_99 vdd gnd cell_6t
Xbit_r100_c62 bl_62 br_62 wl_100 vdd gnd cell_6t
Xbit_r101_c62 bl_62 br_62 wl_101 vdd gnd cell_6t
Xbit_r102_c62 bl_62 br_62 wl_102 vdd gnd cell_6t
Xbit_r103_c62 bl_62 br_62 wl_103 vdd gnd cell_6t
Xbit_r104_c62 bl_62 br_62 wl_104 vdd gnd cell_6t
Xbit_r105_c62 bl_62 br_62 wl_105 vdd gnd cell_6t
Xbit_r106_c62 bl_62 br_62 wl_106 vdd gnd cell_6t
Xbit_r107_c62 bl_62 br_62 wl_107 vdd gnd cell_6t
Xbit_r108_c62 bl_62 br_62 wl_108 vdd gnd cell_6t
Xbit_r109_c62 bl_62 br_62 wl_109 vdd gnd cell_6t
Xbit_r110_c62 bl_62 br_62 wl_110 vdd gnd cell_6t
Xbit_r111_c62 bl_62 br_62 wl_111 vdd gnd cell_6t
Xbit_r112_c62 bl_62 br_62 wl_112 vdd gnd cell_6t
Xbit_r113_c62 bl_62 br_62 wl_113 vdd gnd cell_6t
Xbit_r114_c62 bl_62 br_62 wl_114 vdd gnd cell_6t
Xbit_r115_c62 bl_62 br_62 wl_115 vdd gnd cell_6t
Xbit_r116_c62 bl_62 br_62 wl_116 vdd gnd cell_6t
Xbit_r117_c62 bl_62 br_62 wl_117 vdd gnd cell_6t
Xbit_r118_c62 bl_62 br_62 wl_118 vdd gnd cell_6t
Xbit_r119_c62 bl_62 br_62 wl_119 vdd gnd cell_6t
Xbit_r120_c62 bl_62 br_62 wl_120 vdd gnd cell_6t
Xbit_r121_c62 bl_62 br_62 wl_121 vdd gnd cell_6t
Xbit_r122_c62 bl_62 br_62 wl_122 vdd gnd cell_6t
Xbit_r123_c62 bl_62 br_62 wl_123 vdd gnd cell_6t
Xbit_r124_c62 bl_62 br_62 wl_124 vdd gnd cell_6t
Xbit_r125_c62 bl_62 br_62 wl_125 vdd gnd cell_6t
Xbit_r126_c62 bl_62 br_62 wl_126 vdd gnd cell_6t
Xbit_r127_c62 bl_62 br_62 wl_127 vdd gnd cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd cell_6t
Xbit_r1_c63 bl_63 br_63 wl_1 vdd gnd cell_6t
Xbit_r2_c63 bl_63 br_63 wl_2 vdd gnd cell_6t
Xbit_r3_c63 bl_63 br_63 wl_3 vdd gnd cell_6t
Xbit_r4_c63 bl_63 br_63 wl_4 vdd gnd cell_6t
Xbit_r5_c63 bl_63 br_63 wl_5 vdd gnd cell_6t
Xbit_r6_c63 bl_63 br_63 wl_6 vdd gnd cell_6t
Xbit_r7_c63 bl_63 br_63 wl_7 vdd gnd cell_6t
Xbit_r8_c63 bl_63 br_63 wl_8 vdd gnd cell_6t
Xbit_r9_c63 bl_63 br_63 wl_9 vdd gnd cell_6t
Xbit_r10_c63 bl_63 br_63 wl_10 vdd gnd cell_6t
Xbit_r11_c63 bl_63 br_63 wl_11 vdd gnd cell_6t
Xbit_r12_c63 bl_63 br_63 wl_12 vdd gnd cell_6t
Xbit_r13_c63 bl_63 br_63 wl_13 vdd gnd cell_6t
Xbit_r14_c63 bl_63 br_63 wl_14 vdd gnd cell_6t
Xbit_r15_c63 bl_63 br_63 wl_15 vdd gnd cell_6t
Xbit_r16_c63 bl_63 br_63 wl_16 vdd gnd cell_6t
Xbit_r17_c63 bl_63 br_63 wl_17 vdd gnd cell_6t
Xbit_r18_c63 bl_63 br_63 wl_18 vdd gnd cell_6t
Xbit_r19_c63 bl_63 br_63 wl_19 vdd gnd cell_6t
Xbit_r20_c63 bl_63 br_63 wl_20 vdd gnd cell_6t
Xbit_r21_c63 bl_63 br_63 wl_21 vdd gnd cell_6t
Xbit_r22_c63 bl_63 br_63 wl_22 vdd gnd cell_6t
Xbit_r23_c63 bl_63 br_63 wl_23 vdd gnd cell_6t
Xbit_r24_c63 bl_63 br_63 wl_24 vdd gnd cell_6t
Xbit_r25_c63 bl_63 br_63 wl_25 vdd gnd cell_6t
Xbit_r26_c63 bl_63 br_63 wl_26 vdd gnd cell_6t
Xbit_r27_c63 bl_63 br_63 wl_27 vdd gnd cell_6t
Xbit_r28_c63 bl_63 br_63 wl_28 vdd gnd cell_6t
Xbit_r29_c63 bl_63 br_63 wl_29 vdd gnd cell_6t
Xbit_r30_c63 bl_63 br_63 wl_30 vdd gnd cell_6t
Xbit_r31_c63 bl_63 br_63 wl_31 vdd gnd cell_6t
Xbit_r32_c63 bl_63 br_63 wl_32 vdd gnd cell_6t
Xbit_r33_c63 bl_63 br_63 wl_33 vdd gnd cell_6t
Xbit_r34_c63 bl_63 br_63 wl_34 vdd gnd cell_6t
Xbit_r35_c63 bl_63 br_63 wl_35 vdd gnd cell_6t
Xbit_r36_c63 bl_63 br_63 wl_36 vdd gnd cell_6t
Xbit_r37_c63 bl_63 br_63 wl_37 vdd gnd cell_6t
Xbit_r38_c63 bl_63 br_63 wl_38 vdd gnd cell_6t
Xbit_r39_c63 bl_63 br_63 wl_39 vdd gnd cell_6t
Xbit_r40_c63 bl_63 br_63 wl_40 vdd gnd cell_6t
Xbit_r41_c63 bl_63 br_63 wl_41 vdd gnd cell_6t
Xbit_r42_c63 bl_63 br_63 wl_42 vdd gnd cell_6t
Xbit_r43_c63 bl_63 br_63 wl_43 vdd gnd cell_6t
Xbit_r44_c63 bl_63 br_63 wl_44 vdd gnd cell_6t
Xbit_r45_c63 bl_63 br_63 wl_45 vdd gnd cell_6t
Xbit_r46_c63 bl_63 br_63 wl_46 vdd gnd cell_6t
Xbit_r47_c63 bl_63 br_63 wl_47 vdd gnd cell_6t
Xbit_r48_c63 bl_63 br_63 wl_48 vdd gnd cell_6t
Xbit_r49_c63 bl_63 br_63 wl_49 vdd gnd cell_6t
Xbit_r50_c63 bl_63 br_63 wl_50 vdd gnd cell_6t
Xbit_r51_c63 bl_63 br_63 wl_51 vdd gnd cell_6t
Xbit_r52_c63 bl_63 br_63 wl_52 vdd gnd cell_6t
Xbit_r53_c63 bl_63 br_63 wl_53 vdd gnd cell_6t
Xbit_r54_c63 bl_63 br_63 wl_54 vdd gnd cell_6t
Xbit_r55_c63 bl_63 br_63 wl_55 vdd gnd cell_6t
Xbit_r56_c63 bl_63 br_63 wl_56 vdd gnd cell_6t
Xbit_r57_c63 bl_63 br_63 wl_57 vdd gnd cell_6t
Xbit_r58_c63 bl_63 br_63 wl_58 vdd gnd cell_6t
Xbit_r59_c63 bl_63 br_63 wl_59 vdd gnd cell_6t
Xbit_r60_c63 bl_63 br_63 wl_60 vdd gnd cell_6t
Xbit_r61_c63 bl_63 br_63 wl_61 vdd gnd cell_6t
Xbit_r62_c63 bl_63 br_63 wl_62 vdd gnd cell_6t
Xbit_r63_c63 bl_63 br_63 wl_63 vdd gnd cell_6t
Xbit_r64_c63 bl_63 br_63 wl_64 vdd gnd cell_6t
Xbit_r65_c63 bl_63 br_63 wl_65 vdd gnd cell_6t
Xbit_r66_c63 bl_63 br_63 wl_66 vdd gnd cell_6t
Xbit_r67_c63 bl_63 br_63 wl_67 vdd gnd cell_6t
Xbit_r68_c63 bl_63 br_63 wl_68 vdd gnd cell_6t
Xbit_r69_c63 bl_63 br_63 wl_69 vdd gnd cell_6t
Xbit_r70_c63 bl_63 br_63 wl_70 vdd gnd cell_6t
Xbit_r71_c63 bl_63 br_63 wl_71 vdd gnd cell_6t
Xbit_r72_c63 bl_63 br_63 wl_72 vdd gnd cell_6t
Xbit_r73_c63 bl_63 br_63 wl_73 vdd gnd cell_6t
Xbit_r74_c63 bl_63 br_63 wl_74 vdd gnd cell_6t
Xbit_r75_c63 bl_63 br_63 wl_75 vdd gnd cell_6t
Xbit_r76_c63 bl_63 br_63 wl_76 vdd gnd cell_6t
Xbit_r77_c63 bl_63 br_63 wl_77 vdd gnd cell_6t
Xbit_r78_c63 bl_63 br_63 wl_78 vdd gnd cell_6t
Xbit_r79_c63 bl_63 br_63 wl_79 vdd gnd cell_6t
Xbit_r80_c63 bl_63 br_63 wl_80 vdd gnd cell_6t
Xbit_r81_c63 bl_63 br_63 wl_81 vdd gnd cell_6t
Xbit_r82_c63 bl_63 br_63 wl_82 vdd gnd cell_6t
Xbit_r83_c63 bl_63 br_63 wl_83 vdd gnd cell_6t
Xbit_r84_c63 bl_63 br_63 wl_84 vdd gnd cell_6t
Xbit_r85_c63 bl_63 br_63 wl_85 vdd gnd cell_6t
Xbit_r86_c63 bl_63 br_63 wl_86 vdd gnd cell_6t
Xbit_r87_c63 bl_63 br_63 wl_87 vdd gnd cell_6t
Xbit_r88_c63 bl_63 br_63 wl_88 vdd gnd cell_6t
Xbit_r89_c63 bl_63 br_63 wl_89 vdd gnd cell_6t
Xbit_r90_c63 bl_63 br_63 wl_90 vdd gnd cell_6t
Xbit_r91_c63 bl_63 br_63 wl_91 vdd gnd cell_6t
Xbit_r92_c63 bl_63 br_63 wl_92 vdd gnd cell_6t
Xbit_r93_c63 bl_63 br_63 wl_93 vdd gnd cell_6t
Xbit_r94_c63 bl_63 br_63 wl_94 vdd gnd cell_6t
Xbit_r95_c63 bl_63 br_63 wl_95 vdd gnd cell_6t
Xbit_r96_c63 bl_63 br_63 wl_96 vdd gnd cell_6t
Xbit_r97_c63 bl_63 br_63 wl_97 vdd gnd cell_6t
Xbit_r98_c63 bl_63 br_63 wl_98 vdd gnd cell_6t
Xbit_r99_c63 bl_63 br_63 wl_99 vdd gnd cell_6t
Xbit_r100_c63 bl_63 br_63 wl_100 vdd gnd cell_6t
Xbit_r101_c63 bl_63 br_63 wl_101 vdd gnd cell_6t
Xbit_r102_c63 bl_63 br_63 wl_102 vdd gnd cell_6t
Xbit_r103_c63 bl_63 br_63 wl_103 vdd gnd cell_6t
Xbit_r104_c63 bl_63 br_63 wl_104 vdd gnd cell_6t
Xbit_r105_c63 bl_63 br_63 wl_105 vdd gnd cell_6t
Xbit_r106_c63 bl_63 br_63 wl_106 vdd gnd cell_6t
Xbit_r107_c63 bl_63 br_63 wl_107 vdd gnd cell_6t
Xbit_r108_c63 bl_63 br_63 wl_108 vdd gnd cell_6t
Xbit_r109_c63 bl_63 br_63 wl_109 vdd gnd cell_6t
Xbit_r110_c63 bl_63 br_63 wl_110 vdd gnd cell_6t
Xbit_r111_c63 bl_63 br_63 wl_111 vdd gnd cell_6t
Xbit_r112_c63 bl_63 br_63 wl_112 vdd gnd cell_6t
Xbit_r113_c63 bl_63 br_63 wl_113 vdd gnd cell_6t
Xbit_r114_c63 bl_63 br_63 wl_114 vdd gnd cell_6t
Xbit_r115_c63 bl_63 br_63 wl_115 vdd gnd cell_6t
Xbit_r116_c63 bl_63 br_63 wl_116 vdd gnd cell_6t
Xbit_r117_c63 bl_63 br_63 wl_117 vdd gnd cell_6t
Xbit_r118_c63 bl_63 br_63 wl_118 vdd gnd cell_6t
Xbit_r119_c63 bl_63 br_63 wl_119 vdd gnd cell_6t
Xbit_r120_c63 bl_63 br_63 wl_120 vdd gnd cell_6t
Xbit_r121_c63 bl_63 br_63 wl_121 vdd gnd cell_6t
Xbit_r122_c63 bl_63 br_63 wl_122 vdd gnd cell_6t
Xbit_r123_c63 bl_63 br_63 wl_123 vdd gnd cell_6t
Xbit_r124_c63 bl_63 br_63 wl_124 vdd gnd cell_6t
Xbit_r125_c63 bl_63 br_63 wl_125 vdd gnd cell_6t
Xbit_r126_c63 bl_63 br_63 wl_126 vdd gnd cell_6t
Xbit_r127_c63 bl_63 br_63 wl_127 vdd gnd cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd cell_6t
Xbit_r1_c64 bl_64 br_64 wl_1 vdd gnd cell_6t
Xbit_r2_c64 bl_64 br_64 wl_2 vdd gnd cell_6t
Xbit_r3_c64 bl_64 br_64 wl_3 vdd gnd cell_6t
Xbit_r4_c64 bl_64 br_64 wl_4 vdd gnd cell_6t
Xbit_r5_c64 bl_64 br_64 wl_5 vdd gnd cell_6t
Xbit_r6_c64 bl_64 br_64 wl_6 vdd gnd cell_6t
Xbit_r7_c64 bl_64 br_64 wl_7 vdd gnd cell_6t
Xbit_r8_c64 bl_64 br_64 wl_8 vdd gnd cell_6t
Xbit_r9_c64 bl_64 br_64 wl_9 vdd gnd cell_6t
Xbit_r10_c64 bl_64 br_64 wl_10 vdd gnd cell_6t
Xbit_r11_c64 bl_64 br_64 wl_11 vdd gnd cell_6t
Xbit_r12_c64 bl_64 br_64 wl_12 vdd gnd cell_6t
Xbit_r13_c64 bl_64 br_64 wl_13 vdd gnd cell_6t
Xbit_r14_c64 bl_64 br_64 wl_14 vdd gnd cell_6t
Xbit_r15_c64 bl_64 br_64 wl_15 vdd gnd cell_6t
Xbit_r16_c64 bl_64 br_64 wl_16 vdd gnd cell_6t
Xbit_r17_c64 bl_64 br_64 wl_17 vdd gnd cell_6t
Xbit_r18_c64 bl_64 br_64 wl_18 vdd gnd cell_6t
Xbit_r19_c64 bl_64 br_64 wl_19 vdd gnd cell_6t
Xbit_r20_c64 bl_64 br_64 wl_20 vdd gnd cell_6t
Xbit_r21_c64 bl_64 br_64 wl_21 vdd gnd cell_6t
Xbit_r22_c64 bl_64 br_64 wl_22 vdd gnd cell_6t
Xbit_r23_c64 bl_64 br_64 wl_23 vdd gnd cell_6t
Xbit_r24_c64 bl_64 br_64 wl_24 vdd gnd cell_6t
Xbit_r25_c64 bl_64 br_64 wl_25 vdd gnd cell_6t
Xbit_r26_c64 bl_64 br_64 wl_26 vdd gnd cell_6t
Xbit_r27_c64 bl_64 br_64 wl_27 vdd gnd cell_6t
Xbit_r28_c64 bl_64 br_64 wl_28 vdd gnd cell_6t
Xbit_r29_c64 bl_64 br_64 wl_29 vdd gnd cell_6t
Xbit_r30_c64 bl_64 br_64 wl_30 vdd gnd cell_6t
Xbit_r31_c64 bl_64 br_64 wl_31 vdd gnd cell_6t
Xbit_r32_c64 bl_64 br_64 wl_32 vdd gnd cell_6t
Xbit_r33_c64 bl_64 br_64 wl_33 vdd gnd cell_6t
Xbit_r34_c64 bl_64 br_64 wl_34 vdd gnd cell_6t
Xbit_r35_c64 bl_64 br_64 wl_35 vdd gnd cell_6t
Xbit_r36_c64 bl_64 br_64 wl_36 vdd gnd cell_6t
Xbit_r37_c64 bl_64 br_64 wl_37 vdd gnd cell_6t
Xbit_r38_c64 bl_64 br_64 wl_38 vdd gnd cell_6t
Xbit_r39_c64 bl_64 br_64 wl_39 vdd gnd cell_6t
Xbit_r40_c64 bl_64 br_64 wl_40 vdd gnd cell_6t
Xbit_r41_c64 bl_64 br_64 wl_41 vdd gnd cell_6t
Xbit_r42_c64 bl_64 br_64 wl_42 vdd gnd cell_6t
Xbit_r43_c64 bl_64 br_64 wl_43 vdd gnd cell_6t
Xbit_r44_c64 bl_64 br_64 wl_44 vdd gnd cell_6t
Xbit_r45_c64 bl_64 br_64 wl_45 vdd gnd cell_6t
Xbit_r46_c64 bl_64 br_64 wl_46 vdd gnd cell_6t
Xbit_r47_c64 bl_64 br_64 wl_47 vdd gnd cell_6t
Xbit_r48_c64 bl_64 br_64 wl_48 vdd gnd cell_6t
Xbit_r49_c64 bl_64 br_64 wl_49 vdd gnd cell_6t
Xbit_r50_c64 bl_64 br_64 wl_50 vdd gnd cell_6t
Xbit_r51_c64 bl_64 br_64 wl_51 vdd gnd cell_6t
Xbit_r52_c64 bl_64 br_64 wl_52 vdd gnd cell_6t
Xbit_r53_c64 bl_64 br_64 wl_53 vdd gnd cell_6t
Xbit_r54_c64 bl_64 br_64 wl_54 vdd gnd cell_6t
Xbit_r55_c64 bl_64 br_64 wl_55 vdd gnd cell_6t
Xbit_r56_c64 bl_64 br_64 wl_56 vdd gnd cell_6t
Xbit_r57_c64 bl_64 br_64 wl_57 vdd gnd cell_6t
Xbit_r58_c64 bl_64 br_64 wl_58 vdd gnd cell_6t
Xbit_r59_c64 bl_64 br_64 wl_59 vdd gnd cell_6t
Xbit_r60_c64 bl_64 br_64 wl_60 vdd gnd cell_6t
Xbit_r61_c64 bl_64 br_64 wl_61 vdd gnd cell_6t
Xbit_r62_c64 bl_64 br_64 wl_62 vdd gnd cell_6t
Xbit_r63_c64 bl_64 br_64 wl_63 vdd gnd cell_6t
Xbit_r64_c64 bl_64 br_64 wl_64 vdd gnd cell_6t
Xbit_r65_c64 bl_64 br_64 wl_65 vdd gnd cell_6t
Xbit_r66_c64 bl_64 br_64 wl_66 vdd gnd cell_6t
Xbit_r67_c64 bl_64 br_64 wl_67 vdd gnd cell_6t
Xbit_r68_c64 bl_64 br_64 wl_68 vdd gnd cell_6t
Xbit_r69_c64 bl_64 br_64 wl_69 vdd gnd cell_6t
Xbit_r70_c64 bl_64 br_64 wl_70 vdd gnd cell_6t
Xbit_r71_c64 bl_64 br_64 wl_71 vdd gnd cell_6t
Xbit_r72_c64 bl_64 br_64 wl_72 vdd gnd cell_6t
Xbit_r73_c64 bl_64 br_64 wl_73 vdd gnd cell_6t
Xbit_r74_c64 bl_64 br_64 wl_74 vdd gnd cell_6t
Xbit_r75_c64 bl_64 br_64 wl_75 vdd gnd cell_6t
Xbit_r76_c64 bl_64 br_64 wl_76 vdd gnd cell_6t
Xbit_r77_c64 bl_64 br_64 wl_77 vdd gnd cell_6t
Xbit_r78_c64 bl_64 br_64 wl_78 vdd gnd cell_6t
Xbit_r79_c64 bl_64 br_64 wl_79 vdd gnd cell_6t
Xbit_r80_c64 bl_64 br_64 wl_80 vdd gnd cell_6t
Xbit_r81_c64 bl_64 br_64 wl_81 vdd gnd cell_6t
Xbit_r82_c64 bl_64 br_64 wl_82 vdd gnd cell_6t
Xbit_r83_c64 bl_64 br_64 wl_83 vdd gnd cell_6t
Xbit_r84_c64 bl_64 br_64 wl_84 vdd gnd cell_6t
Xbit_r85_c64 bl_64 br_64 wl_85 vdd gnd cell_6t
Xbit_r86_c64 bl_64 br_64 wl_86 vdd gnd cell_6t
Xbit_r87_c64 bl_64 br_64 wl_87 vdd gnd cell_6t
Xbit_r88_c64 bl_64 br_64 wl_88 vdd gnd cell_6t
Xbit_r89_c64 bl_64 br_64 wl_89 vdd gnd cell_6t
Xbit_r90_c64 bl_64 br_64 wl_90 vdd gnd cell_6t
Xbit_r91_c64 bl_64 br_64 wl_91 vdd gnd cell_6t
Xbit_r92_c64 bl_64 br_64 wl_92 vdd gnd cell_6t
Xbit_r93_c64 bl_64 br_64 wl_93 vdd gnd cell_6t
Xbit_r94_c64 bl_64 br_64 wl_94 vdd gnd cell_6t
Xbit_r95_c64 bl_64 br_64 wl_95 vdd gnd cell_6t
Xbit_r96_c64 bl_64 br_64 wl_96 vdd gnd cell_6t
Xbit_r97_c64 bl_64 br_64 wl_97 vdd gnd cell_6t
Xbit_r98_c64 bl_64 br_64 wl_98 vdd gnd cell_6t
Xbit_r99_c64 bl_64 br_64 wl_99 vdd gnd cell_6t
Xbit_r100_c64 bl_64 br_64 wl_100 vdd gnd cell_6t
Xbit_r101_c64 bl_64 br_64 wl_101 vdd gnd cell_6t
Xbit_r102_c64 bl_64 br_64 wl_102 vdd gnd cell_6t
Xbit_r103_c64 bl_64 br_64 wl_103 vdd gnd cell_6t
Xbit_r104_c64 bl_64 br_64 wl_104 vdd gnd cell_6t
Xbit_r105_c64 bl_64 br_64 wl_105 vdd gnd cell_6t
Xbit_r106_c64 bl_64 br_64 wl_106 vdd gnd cell_6t
Xbit_r107_c64 bl_64 br_64 wl_107 vdd gnd cell_6t
Xbit_r108_c64 bl_64 br_64 wl_108 vdd gnd cell_6t
Xbit_r109_c64 bl_64 br_64 wl_109 vdd gnd cell_6t
Xbit_r110_c64 bl_64 br_64 wl_110 vdd gnd cell_6t
Xbit_r111_c64 bl_64 br_64 wl_111 vdd gnd cell_6t
Xbit_r112_c64 bl_64 br_64 wl_112 vdd gnd cell_6t
Xbit_r113_c64 bl_64 br_64 wl_113 vdd gnd cell_6t
Xbit_r114_c64 bl_64 br_64 wl_114 vdd gnd cell_6t
Xbit_r115_c64 bl_64 br_64 wl_115 vdd gnd cell_6t
Xbit_r116_c64 bl_64 br_64 wl_116 vdd gnd cell_6t
Xbit_r117_c64 bl_64 br_64 wl_117 vdd gnd cell_6t
Xbit_r118_c64 bl_64 br_64 wl_118 vdd gnd cell_6t
Xbit_r119_c64 bl_64 br_64 wl_119 vdd gnd cell_6t
Xbit_r120_c64 bl_64 br_64 wl_120 vdd gnd cell_6t
Xbit_r121_c64 bl_64 br_64 wl_121 vdd gnd cell_6t
Xbit_r122_c64 bl_64 br_64 wl_122 vdd gnd cell_6t
Xbit_r123_c64 bl_64 br_64 wl_123 vdd gnd cell_6t
Xbit_r124_c64 bl_64 br_64 wl_124 vdd gnd cell_6t
Xbit_r125_c64 bl_64 br_64 wl_125 vdd gnd cell_6t
Xbit_r126_c64 bl_64 br_64 wl_126 vdd gnd cell_6t
Xbit_r127_c64 bl_64 br_64 wl_127 vdd gnd cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd cell_6t
Xbit_r1_c65 bl_65 br_65 wl_1 vdd gnd cell_6t
Xbit_r2_c65 bl_65 br_65 wl_2 vdd gnd cell_6t
Xbit_r3_c65 bl_65 br_65 wl_3 vdd gnd cell_6t
Xbit_r4_c65 bl_65 br_65 wl_4 vdd gnd cell_6t
Xbit_r5_c65 bl_65 br_65 wl_5 vdd gnd cell_6t
Xbit_r6_c65 bl_65 br_65 wl_6 vdd gnd cell_6t
Xbit_r7_c65 bl_65 br_65 wl_7 vdd gnd cell_6t
Xbit_r8_c65 bl_65 br_65 wl_8 vdd gnd cell_6t
Xbit_r9_c65 bl_65 br_65 wl_9 vdd gnd cell_6t
Xbit_r10_c65 bl_65 br_65 wl_10 vdd gnd cell_6t
Xbit_r11_c65 bl_65 br_65 wl_11 vdd gnd cell_6t
Xbit_r12_c65 bl_65 br_65 wl_12 vdd gnd cell_6t
Xbit_r13_c65 bl_65 br_65 wl_13 vdd gnd cell_6t
Xbit_r14_c65 bl_65 br_65 wl_14 vdd gnd cell_6t
Xbit_r15_c65 bl_65 br_65 wl_15 vdd gnd cell_6t
Xbit_r16_c65 bl_65 br_65 wl_16 vdd gnd cell_6t
Xbit_r17_c65 bl_65 br_65 wl_17 vdd gnd cell_6t
Xbit_r18_c65 bl_65 br_65 wl_18 vdd gnd cell_6t
Xbit_r19_c65 bl_65 br_65 wl_19 vdd gnd cell_6t
Xbit_r20_c65 bl_65 br_65 wl_20 vdd gnd cell_6t
Xbit_r21_c65 bl_65 br_65 wl_21 vdd gnd cell_6t
Xbit_r22_c65 bl_65 br_65 wl_22 vdd gnd cell_6t
Xbit_r23_c65 bl_65 br_65 wl_23 vdd gnd cell_6t
Xbit_r24_c65 bl_65 br_65 wl_24 vdd gnd cell_6t
Xbit_r25_c65 bl_65 br_65 wl_25 vdd gnd cell_6t
Xbit_r26_c65 bl_65 br_65 wl_26 vdd gnd cell_6t
Xbit_r27_c65 bl_65 br_65 wl_27 vdd gnd cell_6t
Xbit_r28_c65 bl_65 br_65 wl_28 vdd gnd cell_6t
Xbit_r29_c65 bl_65 br_65 wl_29 vdd gnd cell_6t
Xbit_r30_c65 bl_65 br_65 wl_30 vdd gnd cell_6t
Xbit_r31_c65 bl_65 br_65 wl_31 vdd gnd cell_6t
Xbit_r32_c65 bl_65 br_65 wl_32 vdd gnd cell_6t
Xbit_r33_c65 bl_65 br_65 wl_33 vdd gnd cell_6t
Xbit_r34_c65 bl_65 br_65 wl_34 vdd gnd cell_6t
Xbit_r35_c65 bl_65 br_65 wl_35 vdd gnd cell_6t
Xbit_r36_c65 bl_65 br_65 wl_36 vdd gnd cell_6t
Xbit_r37_c65 bl_65 br_65 wl_37 vdd gnd cell_6t
Xbit_r38_c65 bl_65 br_65 wl_38 vdd gnd cell_6t
Xbit_r39_c65 bl_65 br_65 wl_39 vdd gnd cell_6t
Xbit_r40_c65 bl_65 br_65 wl_40 vdd gnd cell_6t
Xbit_r41_c65 bl_65 br_65 wl_41 vdd gnd cell_6t
Xbit_r42_c65 bl_65 br_65 wl_42 vdd gnd cell_6t
Xbit_r43_c65 bl_65 br_65 wl_43 vdd gnd cell_6t
Xbit_r44_c65 bl_65 br_65 wl_44 vdd gnd cell_6t
Xbit_r45_c65 bl_65 br_65 wl_45 vdd gnd cell_6t
Xbit_r46_c65 bl_65 br_65 wl_46 vdd gnd cell_6t
Xbit_r47_c65 bl_65 br_65 wl_47 vdd gnd cell_6t
Xbit_r48_c65 bl_65 br_65 wl_48 vdd gnd cell_6t
Xbit_r49_c65 bl_65 br_65 wl_49 vdd gnd cell_6t
Xbit_r50_c65 bl_65 br_65 wl_50 vdd gnd cell_6t
Xbit_r51_c65 bl_65 br_65 wl_51 vdd gnd cell_6t
Xbit_r52_c65 bl_65 br_65 wl_52 vdd gnd cell_6t
Xbit_r53_c65 bl_65 br_65 wl_53 vdd gnd cell_6t
Xbit_r54_c65 bl_65 br_65 wl_54 vdd gnd cell_6t
Xbit_r55_c65 bl_65 br_65 wl_55 vdd gnd cell_6t
Xbit_r56_c65 bl_65 br_65 wl_56 vdd gnd cell_6t
Xbit_r57_c65 bl_65 br_65 wl_57 vdd gnd cell_6t
Xbit_r58_c65 bl_65 br_65 wl_58 vdd gnd cell_6t
Xbit_r59_c65 bl_65 br_65 wl_59 vdd gnd cell_6t
Xbit_r60_c65 bl_65 br_65 wl_60 vdd gnd cell_6t
Xbit_r61_c65 bl_65 br_65 wl_61 vdd gnd cell_6t
Xbit_r62_c65 bl_65 br_65 wl_62 vdd gnd cell_6t
Xbit_r63_c65 bl_65 br_65 wl_63 vdd gnd cell_6t
Xbit_r64_c65 bl_65 br_65 wl_64 vdd gnd cell_6t
Xbit_r65_c65 bl_65 br_65 wl_65 vdd gnd cell_6t
Xbit_r66_c65 bl_65 br_65 wl_66 vdd gnd cell_6t
Xbit_r67_c65 bl_65 br_65 wl_67 vdd gnd cell_6t
Xbit_r68_c65 bl_65 br_65 wl_68 vdd gnd cell_6t
Xbit_r69_c65 bl_65 br_65 wl_69 vdd gnd cell_6t
Xbit_r70_c65 bl_65 br_65 wl_70 vdd gnd cell_6t
Xbit_r71_c65 bl_65 br_65 wl_71 vdd gnd cell_6t
Xbit_r72_c65 bl_65 br_65 wl_72 vdd gnd cell_6t
Xbit_r73_c65 bl_65 br_65 wl_73 vdd gnd cell_6t
Xbit_r74_c65 bl_65 br_65 wl_74 vdd gnd cell_6t
Xbit_r75_c65 bl_65 br_65 wl_75 vdd gnd cell_6t
Xbit_r76_c65 bl_65 br_65 wl_76 vdd gnd cell_6t
Xbit_r77_c65 bl_65 br_65 wl_77 vdd gnd cell_6t
Xbit_r78_c65 bl_65 br_65 wl_78 vdd gnd cell_6t
Xbit_r79_c65 bl_65 br_65 wl_79 vdd gnd cell_6t
Xbit_r80_c65 bl_65 br_65 wl_80 vdd gnd cell_6t
Xbit_r81_c65 bl_65 br_65 wl_81 vdd gnd cell_6t
Xbit_r82_c65 bl_65 br_65 wl_82 vdd gnd cell_6t
Xbit_r83_c65 bl_65 br_65 wl_83 vdd gnd cell_6t
Xbit_r84_c65 bl_65 br_65 wl_84 vdd gnd cell_6t
Xbit_r85_c65 bl_65 br_65 wl_85 vdd gnd cell_6t
Xbit_r86_c65 bl_65 br_65 wl_86 vdd gnd cell_6t
Xbit_r87_c65 bl_65 br_65 wl_87 vdd gnd cell_6t
Xbit_r88_c65 bl_65 br_65 wl_88 vdd gnd cell_6t
Xbit_r89_c65 bl_65 br_65 wl_89 vdd gnd cell_6t
Xbit_r90_c65 bl_65 br_65 wl_90 vdd gnd cell_6t
Xbit_r91_c65 bl_65 br_65 wl_91 vdd gnd cell_6t
Xbit_r92_c65 bl_65 br_65 wl_92 vdd gnd cell_6t
Xbit_r93_c65 bl_65 br_65 wl_93 vdd gnd cell_6t
Xbit_r94_c65 bl_65 br_65 wl_94 vdd gnd cell_6t
Xbit_r95_c65 bl_65 br_65 wl_95 vdd gnd cell_6t
Xbit_r96_c65 bl_65 br_65 wl_96 vdd gnd cell_6t
Xbit_r97_c65 bl_65 br_65 wl_97 vdd gnd cell_6t
Xbit_r98_c65 bl_65 br_65 wl_98 vdd gnd cell_6t
Xbit_r99_c65 bl_65 br_65 wl_99 vdd gnd cell_6t
Xbit_r100_c65 bl_65 br_65 wl_100 vdd gnd cell_6t
Xbit_r101_c65 bl_65 br_65 wl_101 vdd gnd cell_6t
Xbit_r102_c65 bl_65 br_65 wl_102 vdd gnd cell_6t
Xbit_r103_c65 bl_65 br_65 wl_103 vdd gnd cell_6t
Xbit_r104_c65 bl_65 br_65 wl_104 vdd gnd cell_6t
Xbit_r105_c65 bl_65 br_65 wl_105 vdd gnd cell_6t
Xbit_r106_c65 bl_65 br_65 wl_106 vdd gnd cell_6t
Xbit_r107_c65 bl_65 br_65 wl_107 vdd gnd cell_6t
Xbit_r108_c65 bl_65 br_65 wl_108 vdd gnd cell_6t
Xbit_r109_c65 bl_65 br_65 wl_109 vdd gnd cell_6t
Xbit_r110_c65 bl_65 br_65 wl_110 vdd gnd cell_6t
Xbit_r111_c65 bl_65 br_65 wl_111 vdd gnd cell_6t
Xbit_r112_c65 bl_65 br_65 wl_112 vdd gnd cell_6t
Xbit_r113_c65 bl_65 br_65 wl_113 vdd gnd cell_6t
Xbit_r114_c65 bl_65 br_65 wl_114 vdd gnd cell_6t
Xbit_r115_c65 bl_65 br_65 wl_115 vdd gnd cell_6t
Xbit_r116_c65 bl_65 br_65 wl_116 vdd gnd cell_6t
Xbit_r117_c65 bl_65 br_65 wl_117 vdd gnd cell_6t
Xbit_r118_c65 bl_65 br_65 wl_118 vdd gnd cell_6t
Xbit_r119_c65 bl_65 br_65 wl_119 vdd gnd cell_6t
Xbit_r120_c65 bl_65 br_65 wl_120 vdd gnd cell_6t
Xbit_r121_c65 bl_65 br_65 wl_121 vdd gnd cell_6t
Xbit_r122_c65 bl_65 br_65 wl_122 vdd gnd cell_6t
Xbit_r123_c65 bl_65 br_65 wl_123 vdd gnd cell_6t
Xbit_r124_c65 bl_65 br_65 wl_124 vdd gnd cell_6t
Xbit_r125_c65 bl_65 br_65 wl_125 vdd gnd cell_6t
Xbit_r126_c65 bl_65 br_65 wl_126 vdd gnd cell_6t
Xbit_r127_c65 bl_65 br_65 wl_127 vdd gnd cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd cell_6t
Xbit_r1_c66 bl_66 br_66 wl_1 vdd gnd cell_6t
Xbit_r2_c66 bl_66 br_66 wl_2 vdd gnd cell_6t
Xbit_r3_c66 bl_66 br_66 wl_3 vdd gnd cell_6t
Xbit_r4_c66 bl_66 br_66 wl_4 vdd gnd cell_6t
Xbit_r5_c66 bl_66 br_66 wl_5 vdd gnd cell_6t
Xbit_r6_c66 bl_66 br_66 wl_6 vdd gnd cell_6t
Xbit_r7_c66 bl_66 br_66 wl_7 vdd gnd cell_6t
Xbit_r8_c66 bl_66 br_66 wl_8 vdd gnd cell_6t
Xbit_r9_c66 bl_66 br_66 wl_9 vdd gnd cell_6t
Xbit_r10_c66 bl_66 br_66 wl_10 vdd gnd cell_6t
Xbit_r11_c66 bl_66 br_66 wl_11 vdd gnd cell_6t
Xbit_r12_c66 bl_66 br_66 wl_12 vdd gnd cell_6t
Xbit_r13_c66 bl_66 br_66 wl_13 vdd gnd cell_6t
Xbit_r14_c66 bl_66 br_66 wl_14 vdd gnd cell_6t
Xbit_r15_c66 bl_66 br_66 wl_15 vdd gnd cell_6t
Xbit_r16_c66 bl_66 br_66 wl_16 vdd gnd cell_6t
Xbit_r17_c66 bl_66 br_66 wl_17 vdd gnd cell_6t
Xbit_r18_c66 bl_66 br_66 wl_18 vdd gnd cell_6t
Xbit_r19_c66 bl_66 br_66 wl_19 vdd gnd cell_6t
Xbit_r20_c66 bl_66 br_66 wl_20 vdd gnd cell_6t
Xbit_r21_c66 bl_66 br_66 wl_21 vdd gnd cell_6t
Xbit_r22_c66 bl_66 br_66 wl_22 vdd gnd cell_6t
Xbit_r23_c66 bl_66 br_66 wl_23 vdd gnd cell_6t
Xbit_r24_c66 bl_66 br_66 wl_24 vdd gnd cell_6t
Xbit_r25_c66 bl_66 br_66 wl_25 vdd gnd cell_6t
Xbit_r26_c66 bl_66 br_66 wl_26 vdd gnd cell_6t
Xbit_r27_c66 bl_66 br_66 wl_27 vdd gnd cell_6t
Xbit_r28_c66 bl_66 br_66 wl_28 vdd gnd cell_6t
Xbit_r29_c66 bl_66 br_66 wl_29 vdd gnd cell_6t
Xbit_r30_c66 bl_66 br_66 wl_30 vdd gnd cell_6t
Xbit_r31_c66 bl_66 br_66 wl_31 vdd gnd cell_6t
Xbit_r32_c66 bl_66 br_66 wl_32 vdd gnd cell_6t
Xbit_r33_c66 bl_66 br_66 wl_33 vdd gnd cell_6t
Xbit_r34_c66 bl_66 br_66 wl_34 vdd gnd cell_6t
Xbit_r35_c66 bl_66 br_66 wl_35 vdd gnd cell_6t
Xbit_r36_c66 bl_66 br_66 wl_36 vdd gnd cell_6t
Xbit_r37_c66 bl_66 br_66 wl_37 vdd gnd cell_6t
Xbit_r38_c66 bl_66 br_66 wl_38 vdd gnd cell_6t
Xbit_r39_c66 bl_66 br_66 wl_39 vdd gnd cell_6t
Xbit_r40_c66 bl_66 br_66 wl_40 vdd gnd cell_6t
Xbit_r41_c66 bl_66 br_66 wl_41 vdd gnd cell_6t
Xbit_r42_c66 bl_66 br_66 wl_42 vdd gnd cell_6t
Xbit_r43_c66 bl_66 br_66 wl_43 vdd gnd cell_6t
Xbit_r44_c66 bl_66 br_66 wl_44 vdd gnd cell_6t
Xbit_r45_c66 bl_66 br_66 wl_45 vdd gnd cell_6t
Xbit_r46_c66 bl_66 br_66 wl_46 vdd gnd cell_6t
Xbit_r47_c66 bl_66 br_66 wl_47 vdd gnd cell_6t
Xbit_r48_c66 bl_66 br_66 wl_48 vdd gnd cell_6t
Xbit_r49_c66 bl_66 br_66 wl_49 vdd gnd cell_6t
Xbit_r50_c66 bl_66 br_66 wl_50 vdd gnd cell_6t
Xbit_r51_c66 bl_66 br_66 wl_51 vdd gnd cell_6t
Xbit_r52_c66 bl_66 br_66 wl_52 vdd gnd cell_6t
Xbit_r53_c66 bl_66 br_66 wl_53 vdd gnd cell_6t
Xbit_r54_c66 bl_66 br_66 wl_54 vdd gnd cell_6t
Xbit_r55_c66 bl_66 br_66 wl_55 vdd gnd cell_6t
Xbit_r56_c66 bl_66 br_66 wl_56 vdd gnd cell_6t
Xbit_r57_c66 bl_66 br_66 wl_57 vdd gnd cell_6t
Xbit_r58_c66 bl_66 br_66 wl_58 vdd gnd cell_6t
Xbit_r59_c66 bl_66 br_66 wl_59 vdd gnd cell_6t
Xbit_r60_c66 bl_66 br_66 wl_60 vdd gnd cell_6t
Xbit_r61_c66 bl_66 br_66 wl_61 vdd gnd cell_6t
Xbit_r62_c66 bl_66 br_66 wl_62 vdd gnd cell_6t
Xbit_r63_c66 bl_66 br_66 wl_63 vdd gnd cell_6t
Xbit_r64_c66 bl_66 br_66 wl_64 vdd gnd cell_6t
Xbit_r65_c66 bl_66 br_66 wl_65 vdd gnd cell_6t
Xbit_r66_c66 bl_66 br_66 wl_66 vdd gnd cell_6t
Xbit_r67_c66 bl_66 br_66 wl_67 vdd gnd cell_6t
Xbit_r68_c66 bl_66 br_66 wl_68 vdd gnd cell_6t
Xbit_r69_c66 bl_66 br_66 wl_69 vdd gnd cell_6t
Xbit_r70_c66 bl_66 br_66 wl_70 vdd gnd cell_6t
Xbit_r71_c66 bl_66 br_66 wl_71 vdd gnd cell_6t
Xbit_r72_c66 bl_66 br_66 wl_72 vdd gnd cell_6t
Xbit_r73_c66 bl_66 br_66 wl_73 vdd gnd cell_6t
Xbit_r74_c66 bl_66 br_66 wl_74 vdd gnd cell_6t
Xbit_r75_c66 bl_66 br_66 wl_75 vdd gnd cell_6t
Xbit_r76_c66 bl_66 br_66 wl_76 vdd gnd cell_6t
Xbit_r77_c66 bl_66 br_66 wl_77 vdd gnd cell_6t
Xbit_r78_c66 bl_66 br_66 wl_78 vdd gnd cell_6t
Xbit_r79_c66 bl_66 br_66 wl_79 vdd gnd cell_6t
Xbit_r80_c66 bl_66 br_66 wl_80 vdd gnd cell_6t
Xbit_r81_c66 bl_66 br_66 wl_81 vdd gnd cell_6t
Xbit_r82_c66 bl_66 br_66 wl_82 vdd gnd cell_6t
Xbit_r83_c66 bl_66 br_66 wl_83 vdd gnd cell_6t
Xbit_r84_c66 bl_66 br_66 wl_84 vdd gnd cell_6t
Xbit_r85_c66 bl_66 br_66 wl_85 vdd gnd cell_6t
Xbit_r86_c66 bl_66 br_66 wl_86 vdd gnd cell_6t
Xbit_r87_c66 bl_66 br_66 wl_87 vdd gnd cell_6t
Xbit_r88_c66 bl_66 br_66 wl_88 vdd gnd cell_6t
Xbit_r89_c66 bl_66 br_66 wl_89 vdd gnd cell_6t
Xbit_r90_c66 bl_66 br_66 wl_90 vdd gnd cell_6t
Xbit_r91_c66 bl_66 br_66 wl_91 vdd gnd cell_6t
Xbit_r92_c66 bl_66 br_66 wl_92 vdd gnd cell_6t
Xbit_r93_c66 bl_66 br_66 wl_93 vdd gnd cell_6t
Xbit_r94_c66 bl_66 br_66 wl_94 vdd gnd cell_6t
Xbit_r95_c66 bl_66 br_66 wl_95 vdd gnd cell_6t
Xbit_r96_c66 bl_66 br_66 wl_96 vdd gnd cell_6t
Xbit_r97_c66 bl_66 br_66 wl_97 vdd gnd cell_6t
Xbit_r98_c66 bl_66 br_66 wl_98 vdd gnd cell_6t
Xbit_r99_c66 bl_66 br_66 wl_99 vdd gnd cell_6t
Xbit_r100_c66 bl_66 br_66 wl_100 vdd gnd cell_6t
Xbit_r101_c66 bl_66 br_66 wl_101 vdd gnd cell_6t
Xbit_r102_c66 bl_66 br_66 wl_102 vdd gnd cell_6t
Xbit_r103_c66 bl_66 br_66 wl_103 vdd gnd cell_6t
Xbit_r104_c66 bl_66 br_66 wl_104 vdd gnd cell_6t
Xbit_r105_c66 bl_66 br_66 wl_105 vdd gnd cell_6t
Xbit_r106_c66 bl_66 br_66 wl_106 vdd gnd cell_6t
Xbit_r107_c66 bl_66 br_66 wl_107 vdd gnd cell_6t
Xbit_r108_c66 bl_66 br_66 wl_108 vdd gnd cell_6t
Xbit_r109_c66 bl_66 br_66 wl_109 vdd gnd cell_6t
Xbit_r110_c66 bl_66 br_66 wl_110 vdd gnd cell_6t
Xbit_r111_c66 bl_66 br_66 wl_111 vdd gnd cell_6t
Xbit_r112_c66 bl_66 br_66 wl_112 vdd gnd cell_6t
Xbit_r113_c66 bl_66 br_66 wl_113 vdd gnd cell_6t
Xbit_r114_c66 bl_66 br_66 wl_114 vdd gnd cell_6t
Xbit_r115_c66 bl_66 br_66 wl_115 vdd gnd cell_6t
Xbit_r116_c66 bl_66 br_66 wl_116 vdd gnd cell_6t
Xbit_r117_c66 bl_66 br_66 wl_117 vdd gnd cell_6t
Xbit_r118_c66 bl_66 br_66 wl_118 vdd gnd cell_6t
Xbit_r119_c66 bl_66 br_66 wl_119 vdd gnd cell_6t
Xbit_r120_c66 bl_66 br_66 wl_120 vdd gnd cell_6t
Xbit_r121_c66 bl_66 br_66 wl_121 vdd gnd cell_6t
Xbit_r122_c66 bl_66 br_66 wl_122 vdd gnd cell_6t
Xbit_r123_c66 bl_66 br_66 wl_123 vdd gnd cell_6t
Xbit_r124_c66 bl_66 br_66 wl_124 vdd gnd cell_6t
Xbit_r125_c66 bl_66 br_66 wl_125 vdd gnd cell_6t
Xbit_r126_c66 bl_66 br_66 wl_126 vdd gnd cell_6t
Xbit_r127_c66 bl_66 br_66 wl_127 vdd gnd cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd cell_6t
Xbit_r1_c67 bl_67 br_67 wl_1 vdd gnd cell_6t
Xbit_r2_c67 bl_67 br_67 wl_2 vdd gnd cell_6t
Xbit_r3_c67 bl_67 br_67 wl_3 vdd gnd cell_6t
Xbit_r4_c67 bl_67 br_67 wl_4 vdd gnd cell_6t
Xbit_r5_c67 bl_67 br_67 wl_5 vdd gnd cell_6t
Xbit_r6_c67 bl_67 br_67 wl_6 vdd gnd cell_6t
Xbit_r7_c67 bl_67 br_67 wl_7 vdd gnd cell_6t
Xbit_r8_c67 bl_67 br_67 wl_8 vdd gnd cell_6t
Xbit_r9_c67 bl_67 br_67 wl_9 vdd gnd cell_6t
Xbit_r10_c67 bl_67 br_67 wl_10 vdd gnd cell_6t
Xbit_r11_c67 bl_67 br_67 wl_11 vdd gnd cell_6t
Xbit_r12_c67 bl_67 br_67 wl_12 vdd gnd cell_6t
Xbit_r13_c67 bl_67 br_67 wl_13 vdd gnd cell_6t
Xbit_r14_c67 bl_67 br_67 wl_14 vdd gnd cell_6t
Xbit_r15_c67 bl_67 br_67 wl_15 vdd gnd cell_6t
Xbit_r16_c67 bl_67 br_67 wl_16 vdd gnd cell_6t
Xbit_r17_c67 bl_67 br_67 wl_17 vdd gnd cell_6t
Xbit_r18_c67 bl_67 br_67 wl_18 vdd gnd cell_6t
Xbit_r19_c67 bl_67 br_67 wl_19 vdd gnd cell_6t
Xbit_r20_c67 bl_67 br_67 wl_20 vdd gnd cell_6t
Xbit_r21_c67 bl_67 br_67 wl_21 vdd gnd cell_6t
Xbit_r22_c67 bl_67 br_67 wl_22 vdd gnd cell_6t
Xbit_r23_c67 bl_67 br_67 wl_23 vdd gnd cell_6t
Xbit_r24_c67 bl_67 br_67 wl_24 vdd gnd cell_6t
Xbit_r25_c67 bl_67 br_67 wl_25 vdd gnd cell_6t
Xbit_r26_c67 bl_67 br_67 wl_26 vdd gnd cell_6t
Xbit_r27_c67 bl_67 br_67 wl_27 vdd gnd cell_6t
Xbit_r28_c67 bl_67 br_67 wl_28 vdd gnd cell_6t
Xbit_r29_c67 bl_67 br_67 wl_29 vdd gnd cell_6t
Xbit_r30_c67 bl_67 br_67 wl_30 vdd gnd cell_6t
Xbit_r31_c67 bl_67 br_67 wl_31 vdd gnd cell_6t
Xbit_r32_c67 bl_67 br_67 wl_32 vdd gnd cell_6t
Xbit_r33_c67 bl_67 br_67 wl_33 vdd gnd cell_6t
Xbit_r34_c67 bl_67 br_67 wl_34 vdd gnd cell_6t
Xbit_r35_c67 bl_67 br_67 wl_35 vdd gnd cell_6t
Xbit_r36_c67 bl_67 br_67 wl_36 vdd gnd cell_6t
Xbit_r37_c67 bl_67 br_67 wl_37 vdd gnd cell_6t
Xbit_r38_c67 bl_67 br_67 wl_38 vdd gnd cell_6t
Xbit_r39_c67 bl_67 br_67 wl_39 vdd gnd cell_6t
Xbit_r40_c67 bl_67 br_67 wl_40 vdd gnd cell_6t
Xbit_r41_c67 bl_67 br_67 wl_41 vdd gnd cell_6t
Xbit_r42_c67 bl_67 br_67 wl_42 vdd gnd cell_6t
Xbit_r43_c67 bl_67 br_67 wl_43 vdd gnd cell_6t
Xbit_r44_c67 bl_67 br_67 wl_44 vdd gnd cell_6t
Xbit_r45_c67 bl_67 br_67 wl_45 vdd gnd cell_6t
Xbit_r46_c67 bl_67 br_67 wl_46 vdd gnd cell_6t
Xbit_r47_c67 bl_67 br_67 wl_47 vdd gnd cell_6t
Xbit_r48_c67 bl_67 br_67 wl_48 vdd gnd cell_6t
Xbit_r49_c67 bl_67 br_67 wl_49 vdd gnd cell_6t
Xbit_r50_c67 bl_67 br_67 wl_50 vdd gnd cell_6t
Xbit_r51_c67 bl_67 br_67 wl_51 vdd gnd cell_6t
Xbit_r52_c67 bl_67 br_67 wl_52 vdd gnd cell_6t
Xbit_r53_c67 bl_67 br_67 wl_53 vdd gnd cell_6t
Xbit_r54_c67 bl_67 br_67 wl_54 vdd gnd cell_6t
Xbit_r55_c67 bl_67 br_67 wl_55 vdd gnd cell_6t
Xbit_r56_c67 bl_67 br_67 wl_56 vdd gnd cell_6t
Xbit_r57_c67 bl_67 br_67 wl_57 vdd gnd cell_6t
Xbit_r58_c67 bl_67 br_67 wl_58 vdd gnd cell_6t
Xbit_r59_c67 bl_67 br_67 wl_59 vdd gnd cell_6t
Xbit_r60_c67 bl_67 br_67 wl_60 vdd gnd cell_6t
Xbit_r61_c67 bl_67 br_67 wl_61 vdd gnd cell_6t
Xbit_r62_c67 bl_67 br_67 wl_62 vdd gnd cell_6t
Xbit_r63_c67 bl_67 br_67 wl_63 vdd gnd cell_6t
Xbit_r64_c67 bl_67 br_67 wl_64 vdd gnd cell_6t
Xbit_r65_c67 bl_67 br_67 wl_65 vdd gnd cell_6t
Xbit_r66_c67 bl_67 br_67 wl_66 vdd gnd cell_6t
Xbit_r67_c67 bl_67 br_67 wl_67 vdd gnd cell_6t
Xbit_r68_c67 bl_67 br_67 wl_68 vdd gnd cell_6t
Xbit_r69_c67 bl_67 br_67 wl_69 vdd gnd cell_6t
Xbit_r70_c67 bl_67 br_67 wl_70 vdd gnd cell_6t
Xbit_r71_c67 bl_67 br_67 wl_71 vdd gnd cell_6t
Xbit_r72_c67 bl_67 br_67 wl_72 vdd gnd cell_6t
Xbit_r73_c67 bl_67 br_67 wl_73 vdd gnd cell_6t
Xbit_r74_c67 bl_67 br_67 wl_74 vdd gnd cell_6t
Xbit_r75_c67 bl_67 br_67 wl_75 vdd gnd cell_6t
Xbit_r76_c67 bl_67 br_67 wl_76 vdd gnd cell_6t
Xbit_r77_c67 bl_67 br_67 wl_77 vdd gnd cell_6t
Xbit_r78_c67 bl_67 br_67 wl_78 vdd gnd cell_6t
Xbit_r79_c67 bl_67 br_67 wl_79 vdd gnd cell_6t
Xbit_r80_c67 bl_67 br_67 wl_80 vdd gnd cell_6t
Xbit_r81_c67 bl_67 br_67 wl_81 vdd gnd cell_6t
Xbit_r82_c67 bl_67 br_67 wl_82 vdd gnd cell_6t
Xbit_r83_c67 bl_67 br_67 wl_83 vdd gnd cell_6t
Xbit_r84_c67 bl_67 br_67 wl_84 vdd gnd cell_6t
Xbit_r85_c67 bl_67 br_67 wl_85 vdd gnd cell_6t
Xbit_r86_c67 bl_67 br_67 wl_86 vdd gnd cell_6t
Xbit_r87_c67 bl_67 br_67 wl_87 vdd gnd cell_6t
Xbit_r88_c67 bl_67 br_67 wl_88 vdd gnd cell_6t
Xbit_r89_c67 bl_67 br_67 wl_89 vdd gnd cell_6t
Xbit_r90_c67 bl_67 br_67 wl_90 vdd gnd cell_6t
Xbit_r91_c67 bl_67 br_67 wl_91 vdd gnd cell_6t
Xbit_r92_c67 bl_67 br_67 wl_92 vdd gnd cell_6t
Xbit_r93_c67 bl_67 br_67 wl_93 vdd gnd cell_6t
Xbit_r94_c67 bl_67 br_67 wl_94 vdd gnd cell_6t
Xbit_r95_c67 bl_67 br_67 wl_95 vdd gnd cell_6t
Xbit_r96_c67 bl_67 br_67 wl_96 vdd gnd cell_6t
Xbit_r97_c67 bl_67 br_67 wl_97 vdd gnd cell_6t
Xbit_r98_c67 bl_67 br_67 wl_98 vdd gnd cell_6t
Xbit_r99_c67 bl_67 br_67 wl_99 vdd gnd cell_6t
Xbit_r100_c67 bl_67 br_67 wl_100 vdd gnd cell_6t
Xbit_r101_c67 bl_67 br_67 wl_101 vdd gnd cell_6t
Xbit_r102_c67 bl_67 br_67 wl_102 vdd gnd cell_6t
Xbit_r103_c67 bl_67 br_67 wl_103 vdd gnd cell_6t
Xbit_r104_c67 bl_67 br_67 wl_104 vdd gnd cell_6t
Xbit_r105_c67 bl_67 br_67 wl_105 vdd gnd cell_6t
Xbit_r106_c67 bl_67 br_67 wl_106 vdd gnd cell_6t
Xbit_r107_c67 bl_67 br_67 wl_107 vdd gnd cell_6t
Xbit_r108_c67 bl_67 br_67 wl_108 vdd gnd cell_6t
Xbit_r109_c67 bl_67 br_67 wl_109 vdd gnd cell_6t
Xbit_r110_c67 bl_67 br_67 wl_110 vdd gnd cell_6t
Xbit_r111_c67 bl_67 br_67 wl_111 vdd gnd cell_6t
Xbit_r112_c67 bl_67 br_67 wl_112 vdd gnd cell_6t
Xbit_r113_c67 bl_67 br_67 wl_113 vdd gnd cell_6t
Xbit_r114_c67 bl_67 br_67 wl_114 vdd gnd cell_6t
Xbit_r115_c67 bl_67 br_67 wl_115 vdd gnd cell_6t
Xbit_r116_c67 bl_67 br_67 wl_116 vdd gnd cell_6t
Xbit_r117_c67 bl_67 br_67 wl_117 vdd gnd cell_6t
Xbit_r118_c67 bl_67 br_67 wl_118 vdd gnd cell_6t
Xbit_r119_c67 bl_67 br_67 wl_119 vdd gnd cell_6t
Xbit_r120_c67 bl_67 br_67 wl_120 vdd gnd cell_6t
Xbit_r121_c67 bl_67 br_67 wl_121 vdd gnd cell_6t
Xbit_r122_c67 bl_67 br_67 wl_122 vdd gnd cell_6t
Xbit_r123_c67 bl_67 br_67 wl_123 vdd gnd cell_6t
Xbit_r124_c67 bl_67 br_67 wl_124 vdd gnd cell_6t
Xbit_r125_c67 bl_67 br_67 wl_125 vdd gnd cell_6t
Xbit_r126_c67 bl_67 br_67 wl_126 vdd gnd cell_6t
Xbit_r127_c67 bl_67 br_67 wl_127 vdd gnd cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd cell_6t
Xbit_r1_c68 bl_68 br_68 wl_1 vdd gnd cell_6t
Xbit_r2_c68 bl_68 br_68 wl_2 vdd gnd cell_6t
Xbit_r3_c68 bl_68 br_68 wl_3 vdd gnd cell_6t
Xbit_r4_c68 bl_68 br_68 wl_4 vdd gnd cell_6t
Xbit_r5_c68 bl_68 br_68 wl_5 vdd gnd cell_6t
Xbit_r6_c68 bl_68 br_68 wl_6 vdd gnd cell_6t
Xbit_r7_c68 bl_68 br_68 wl_7 vdd gnd cell_6t
Xbit_r8_c68 bl_68 br_68 wl_8 vdd gnd cell_6t
Xbit_r9_c68 bl_68 br_68 wl_9 vdd gnd cell_6t
Xbit_r10_c68 bl_68 br_68 wl_10 vdd gnd cell_6t
Xbit_r11_c68 bl_68 br_68 wl_11 vdd gnd cell_6t
Xbit_r12_c68 bl_68 br_68 wl_12 vdd gnd cell_6t
Xbit_r13_c68 bl_68 br_68 wl_13 vdd gnd cell_6t
Xbit_r14_c68 bl_68 br_68 wl_14 vdd gnd cell_6t
Xbit_r15_c68 bl_68 br_68 wl_15 vdd gnd cell_6t
Xbit_r16_c68 bl_68 br_68 wl_16 vdd gnd cell_6t
Xbit_r17_c68 bl_68 br_68 wl_17 vdd gnd cell_6t
Xbit_r18_c68 bl_68 br_68 wl_18 vdd gnd cell_6t
Xbit_r19_c68 bl_68 br_68 wl_19 vdd gnd cell_6t
Xbit_r20_c68 bl_68 br_68 wl_20 vdd gnd cell_6t
Xbit_r21_c68 bl_68 br_68 wl_21 vdd gnd cell_6t
Xbit_r22_c68 bl_68 br_68 wl_22 vdd gnd cell_6t
Xbit_r23_c68 bl_68 br_68 wl_23 vdd gnd cell_6t
Xbit_r24_c68 bl_68 br_68 wl_24 vdd gnd cell_6t
Xbit_r25_c68 bl_68 br_68 wl_25 vdd gnd cell_6t
Xbit_r26_c68 bl_68 br_68 wl_26 vdd gnd cell_6t
Xbit_r27_c68 bl_68 br_68 wl_27 vdd gnd cell_6t
Xbit_r28_c68 bl_68 br_68 wl_28 vdd gnd cell_6t
Xbit_r29_c68 bl_68 br_68 wl_29 vdd gnd cell_6t
Xbit_r30_c68 bl_68 br_68 wl_30 vdd gnd cell_6t
Xbit_r31_c68 bl_68 br_68 wl_31 vdd gnd cell_6t
Xbit_r32_c68 bl_68 br_68 wl_32 vdd gnd cell_6t
Xbit_r33_c68 bl_68 br_68 wl_33 vdd gnd cell_6t
Xbit_r34_c68 bl_68 br_68 wl_34 vdd gnd cell_6t
Xbit_r35_c68 bl_68 br_68 wl_35 vdd gnd cell_6t
Xbit_r36_c68 bl_68 br_68 wl_36 vdd gnd cell_6t
Xbit_r37_c68 bl_68 br_68 wl_37 vdd gnd cell_6t
Xbit_r38_c68 bl_68 br_68 wl_38 vdd gnd cell_6t
Xbit_r39_c68 bl_68 br_68 wl_39 vdd gnd cell_6t
Xbit_r40_c68 bl_68 br_68 wl_40 vdd gnd cell_6t
Xbit_r41_c68 bl_68 br_68 wl_41 vdd gnd cell_6t
Xbit_r42_c68 bl_68 br_68 wl_42 vdd gnd cell_6t
Xbit_r43_c68 bl_68 br_68 wl_43 vdd gnd cell_6t
Xbit_r44_c68 bl_68 br_68 wl_44 vdd gnd cell_6t
Xbit_r45_c68 bl_68 br_68 wl_45 vdd gnd cell_6t
Xbit_r46_c68 bl_68 br_68 wl_46 vdd gnd cell_6t
Xbit_r47_c68 bl_68 br_68 wl_47 vdd gnd cell_6t
Xbit_r48_c68 bl_68 br_68 wl_48 vdd gnd cell_6t
Xbit_r49_c68 bl_68 br_68 wl_49 vdd gnd cell_6t
Xbit_r50_c68 bl_68 br_68 wl_50 vdd gnd cell_6t
Xbit_r51_c68 bl_68 br_68 wl_51 vdd gnd cell_6t
Xbit_r52_c68 bl_68 br_68 wl_52 vdd gnd cell_6t
Xbit_r53_c68 bl_68 br_68 wl_53 vdd gnd cell_6t
Xbit_r54_c68 bl_68 br_68 wl_54 vdd gnd cell_6t
Xbit_r55_c68 bl_68 br_68 wl_55 vdd gnd cell_6t
Xbit_r56_c68 bl_68 br_68 wl_56 vdd gnd cell_6t
Xbit_r57_c68 bl_68 br_68 wl_57 vdd gnd cell_6t
Xbit_r58_c68 bl_68 br_68 wl_58 vdd gnd cell_6t
Xbit_r59_c68 bl_68 br_68 wl_59 vdd gnd cell_6t
Xbit_r60_c68 bl_68 br_68 wl_60 vdd gnd cell_6t
Xbit_r61_c68 bl_68 br_68 wl_61 vdd gnd cell_6t
Xbit_r62_c68 bl_68 br_68 wl_62 vdd gnd cell_6t
Xbit_r63_c68 bl_68 br_68 wl_63 vdd gnd cell_6t
Xbit_r64_c68 bl_68 br_68 wl_64 vdd gnd cell_6t
Xbit_r65_c68 bl_68 br_68 wl_65 vdd gnd cell_6t
Xbit_r66_c68 bl_68 br_68 wl_66 vdd gnd cell_6t
Xbit_r67_c68 bl_68 br_68 wl_67 vdd gnd cell_6t
Xbit_r68_c68 bl_68 br_68 wl_68 vdd gnd cell_6t
Xbit_r69_c68 bl_68 br_68 wl_69 vdd gnd cell_6t
Xbit_r70_c68 bl_68 br_68 wl_70 vdd gnd cell_6t
Xbit_r71_c68 bl_68 br_68 wl_71 vdd gnd cell_6t
Xbit_r72_c68 bl_68 br_68 wl_72 vdd gnd cell_6t
Xbit_r73_c68 bl_68 br_68 wl_73 vdd gnd cell_6t
Xbit_r74_c68 bl_68 br_68 wl_74 vdd gnd cell_6t
Xbit_r75_c68 bl_68 br_68 wl_75 vdd gnd cell_6t
Xbit_r76_c68 bl_68 br_68 wl_76 vdd gnd cell_6t
Xbit_r77_c68 bl_68 br_68 wl_77 vdd gnd cell_6t
Xbit_r78_c68 bl_68 br_68 wl_78 vdd gnd cell_6t
Xbit_r79_c68 bl_68 br_68 wl_79 vdd gnd cell_6t
Xbit_r80_c68 bl_68 br_68 wl_80 vdd gnd cell_6t
Xbit_r81_c68 bl_68 br_68 wl_81 vdd gnd cell_6t
Xbit_r82_c68 bl_68 br_68 wl_82 vdd gnd cell_6t
Xbit_r83_c68 bl_68 br_68 wl_83 vdd gnd cell_6t
Xbit_r84_c68 bl_68 br_68 wl_84 vdd gnd cell_6t
Xbit_r85_c68 bl_68 br_68 wl_85 vdd gnd cell_6t
Xbit_r86_c68 bl_68 br_68 wl_86 vdd gnd cell_6t
Xbit_r87_c68 bl_68 br_68 wl_87 vdd gnd cell_6t
Xbit_r88_c68 bl_68 br_68 wl_88 vdd gnd cell_6t
Xbit_r89_c68 bl_68 br_68 wl_89 vdd gnd cell_6t
Xbit_r90_c68 bl_68 br_68 wl_90 vdd gnd cell_6t
Xbit_r91_c68 bl_68 br_68 wl_91 vdd gnd cell_6t
Xbit_r92_c68 bl_68 br_68 wl_92 vdd gnd cell_6t
Xbit_r93_c68 bl_68 br_68 wl_93 vdd gnd cell_6t
Xbit_r94_c68 bl_68 br_68 wl_94 vdd gnd cell_6t
Xbit_r95_c68 bl_68 br_68 wl_95 vdd gnd cell_6t
Xbit_r96_c68 bl_68 br_68 wl_96 vdd gnd cell_6t
Xbit_r97_c68 bl_68 br_68 wl_97 vdd gnd cell_6t
Xbit_r98_c68 bl_68 br_68 wl_98 vdd gnd cell_6t
Xbit_r99_c68 bl_68 br_68 wl_99 vdd gnd cell_6t
Xbit_r100_c68 bl_68 br_68 wl_100 vdd gnd cell_6t
Xbit_r101_c68 bl_68 br_68 wl_101 vdd gnd cell_6t
Xbit_r102_c68 bl_68 br_68 wl_102 vdd gnd cell_6t
Xbit_r103_c68 bl_68 br_68 wl_103 vdd gnd cell_6t
Xbit_r104_c68 bl_68 br_68 wl_104 vdd gnd cell_6t
Xbit_r105_c68 bl_68 br_68 wl_105 vdd gnd cell_6t
Xbit_r106_c68 bl_68 br_68 wl_106 vdd gnd cell_6t
Xbit_r107_c68 bl_68 br_68 wl_107 vdd gnd cell_6t
Xbit_r108_c68 bl_68 br_68 wl_108 vdd gnd cell_6t
Xbit_r109_c68 bl_68 br_68 wl_109 vdd gnd cell_6t
Xbit_r110_c68 bl_68 br_68 wl_110 vdd gnd cell_6t
Xbit_r111_c68 bl_68 br_68 wl_111 vdd gnd cell_6t
Xbit_r112_c68 bl_68 br_68 wl_112 vdd gnd cell_6t
Xbit_r113_c68 bl_68 br_68 wl_113 vdd gnd cell_6t
Xbit_r114_c68 bl_68 br_68 wl_114 vdd gnd cell_6t
Xbit_r115_c68 bl_68 br_68 wl_115 vdd gnd cell_6t
Xbit_r116_c68 bl_68 br_68 wl_116 vdd gnd cell_6t
Xbit_r117_c68 bl_68 br_68 wl_117 vdd gnd cell_6t
Xbit_r118_c68 bl_68 br_68 wl_118 vdd gnd cell_6t
Xbit_r119_c68 bl_68 br_68 wl_119 vdd gnd cell_6t
Xbit_r120_c68 bl_68 br_68 wl_120 vdd gnd cell_6t
Xbit_r121_c68 bl_68 br_68 wl_121 vdd gnd cell_6t
Xbit_r122_c68 bl_68 br_68 wl_122 vdd gnd cell_6t
Xbit_r123_c68 bl_68 br_68 wl_123 vdd gnd cell_6t
Xbit_r124_c68 bl_68 br_68 wl_124 vdd gnd cell_6t
Xbit_r125_c68 bl_68 br_68 wl_125 vdd gnd cell_6t
Xbit_r126_c68 bl_68 br_68 wl_126 vdd gnd cell_6t
Xbit_r127_c68 bl_68 br_68 wl_127 vdd gnd cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd cell_6t
Xbit_r1_c69 bl_69 br_69 wl_1 vdd gnd cell_6t
Xbit_r2_c69 bl_69 br_69 wl_2 vdd gnd cell_6t
Xbit_r3_c69 bl_69 br_69 wl_3 vdd gnd cell_6t
Xbit_r4_c69 bl_69 br_69 wl_4 vdd gnd cell_6t
Xbit_r5_c69 bl_69 br_69 wl_5 vdd gnd cell_6t
Xbit_r6_c69 bl_69 br_69 wl_6 vdd gnd cell_6t
Xbit_r7_c69 bl_69 br_69 wl_7 vdd gnd cell_6t
Xbit_r8_c69 bl_69 br_69 wl_8 vdd gnd cell_6t
Xbit_r9_c69 bl_69 br_69 wl_9 vdd gnd cell_6t
Xbit_r10_c69 bl_69 br_69 wl_10 vdd gnd cell_6t
Xbit_r11_c69 bl_69 br_69 wl_11 vdd gnd cell_6t
Xbit_r12_c69 bl_69 br_69 wl_12 vdd gnd cell_6t
Xbit_r13_c69 bl_69 br_69 wl_13 vdd gnd cell_6t
Xbit_r14_c69 bl_69 br_69 wl_14 vdd gnd cell_6t
Xbit_r15_c69 bl_69 br_69 wl_15 vdd gnd cell_6t
Xbit_r16_c69 bl_69 br_69 wl_16 vdd gnd cell_6t
Xbit_r17_c69 bl_69 br_69 wl_17 vdd gnd cell_6t
Xbit_r18_c69 bl_69 br_69 wl_18 vdd gnd cell_6t
Xbit_r19_c69 bl_69 br_69 wl_19 vdd gnd cell_6t
Xbit_r20_c69 bl_69 br_69 wl_20 vdd gnd cell_6t
Xbit_r21_c69 bl_69 br_69 wl_21 vdd gnd cell_6t
Xbit_r22_c69 bl_69 br_69 wl_22 vdd gnd cell_6t
Xbit_r23_c69 bl_69 br_69 wl_23 vdd gnd cell_6t
Xbit_r24_c69 bl_69 br_69 wl_24 vdd gnd cell_6t
Xbit_r25_c69 bl_69 br_69 wl_25 vdd gnd cell_6t
Xbit_r26_c69 bl_69 br_69 wl_26 vdd gnd cell_6t
Xbit_r27_c69 bl_69 br_69 wl_27 vdd gnd cell_6t
Xbit_r28_c69 bl_69 br_69 wl_28 vdd gnd cell_6t
Xbit_r29_c69 bl_69 br_69 wl_29 vdd gnd cell_6t
Xbit_r30_c69 bl_69 br_69 wl_30 vdd gnd cell_6t
Xbit_r31_c69 bl_69 br_69 wl_31 vdd gnd cell_6t
Xbit_r32_c69 bl_69 br_69 wl_32 vdd gnd cell_6t
Xbit_r33_c69 bl_69 br_69 wl_33 vdd gnd cell_6t
Xbit_r34_c69 bl_69 br_69 wl_34 vdd gnd cell_6t
Xbit_r35_c69 bl_69 br_69 wl_35 vdd gnd cell_6t
Xbit_r36_c69 bl_69 br_69 wl_36 vdd gnd cell_6t
Xbit_r37_c69 bl_69 br_69 wl_37 vdd gnd cell_6t
Xbit_r38_c69 bl_69 br_69 wl_38 vdd gnd cell_6t
Xbit_r39_c69 bl_69 br_69 wl_39 vdd gnd cell_6t
Xbit_r40_c69 bl_69 br_69 wl_40 vdd gnd cell_6t
Xbit_r41_c69 bl_69 br_69 wl_41 vdd gnd cell_6t
Xbit_r42_c69 bl_69 br_69 wl_42 vdd gnd cell_6t
Xbit_r43_c69 bl_69 br_69 wl_43 vdd gnd cell_6t
Xbit_r44_c69 bl_69 br_69 wl_44 vdd gnd cell_6t
Xbit_r45_c69 bl_69 br_69 wl_45 vdd gnd cell_6t
Xbit_r46_c69 bl_69 br_69 wl_46 vdd gnd cell_6t
Xbit_r47_c69 bl_69 br_69 wl_47 vdd gnd cell_6t
Xbit_r48_c69 bl_69 br_69 wl_48 vdd gnd cell_6t
Xbit_r49_c69 bl_69 br_69 wl_49 vdd gnd cell_6t
Xbit_r50_c69 bl_69 br_69 wl_50 vdd gnd cell_6t
Xbit_r51_c69 bl_69 br_69 wl_51 vdd gnd cell_6t
Xbit_r52_c69 bl_69 br_69 wl_52 vdd gnd cell_6t
Xbit_r53_c69 bl_69 br_69 wl_53 vdd gnd cell_6t
Xbit_r54_c69 bl_69 br_69 wl_54 vdd gnd cell_6t
Xbit_r55_c69 bl_69 br_69 wl_55 vdd gnd cell_6t
Xbit_r56_c69 bl_69 br_69 wl_56 vdd gnd cell_6t
Xbit_r57_c69 bl_69 br_69 wl_57 vdd gnd cell_6t
Xbit_r58_c69 bl_69 br_69 wl_58 vdd gnd cell_6t
Xbit_r59_c69 bl_69 br_69 wl_59 vdd gnd cell_6t
Xbit_r60_c69 bl_69 br_69 wl_60 vdd gnd cell_6t
Xbit_r61_c69 bl_69 br_69 wl_61 vdd gnd cell_6t
Xbit_r62_c69 bl_69 br_69 wl_62 vdd gnd cell_6t
Xbit_r63_c69 bl_69 br_69 wl_63 vdd gnd cell_6t
Xbit_r64_c69 bl_69 br_69 wl_64 vdd gnd cell_6t
Xbit_r65_c69 bl_69 br_69 wl_65 vdd gnd cell_6t
Xbit_r66_c69 bl_69 br_69 wl_66 vdd gnd cell_6t
Xbit_r67_c69 bl_69 br_69 wl_67 vdd gnd cell_6t
Xbit_r68_c69 bl_69 br_69 wl_68 vdd gnd cell_6t
Xbit_r69_c69 bl_69 br_69 wl_69 vdd gnd cell_6t
Xbit_r70_c69 bl_69 br_69 wl_70 vdd gnd cell_6t
Xbit_r71_c69 bl_69 br_69 wl_71 vdd gnd cell_6t
Xbit_r72_c69 bl_69 br_69 wl_72 vdd gnd cell_6t
Xbit_r73_c69 bl_69 br_69 wl_73 vdd gnd cell_6t
Xbit_r74_c69 bl_69 br_69 wl_74 vdd gnd cell_6t
Xbit_r75_c69 bl_69 br_69 wl_75 vdd gnd cell_6t
Xbit_r76_c69 bl_69 br_69 wl_76 vdd gnd cell_6t
Xbit_r77_c69 bl_69 br_69 wl_77 vdd gnd cell_6t
Xbit_r78_c69 bl_69 br_69 wl_78 vdd gnd cell_6t
Xbit_r79_c69 bl_69 br_69 wl_79 vdd gnd cell_6t
Xbit_r80_c69 bl_69 br_69 wl_80 vdd gnd cell_6t
Xbit_r81_c69 bl_69 br_69 wl_81 vdd gnd cell_6t
Xbit_r82_c69 bl_69 br_69 wl_82 vdd gnd cell_6t
Xbit_r83_c69 bl_69 br_69 wl_83 vdd gnd cell_6t
Xbit_r84_c69 bl_69 br_69 wl_84 vdd gnd cell_6t
Xbit_r85_c69 bl_69 br_69 wl_85 vdd gnd cell_6t
Xbit_r86_c69 bl_69 br_69 wl_86 vdd gnd cell_6t
Xbit_r87_c69 bl_69 br_69 wl_87 vdd gnd cell_6t
Xbit_r88_c69 bl_69 br_69 wl_88 vdd gnd cell_6t
Xbit_r89_c69 bl_69 br_69 wl_89 vdd gnd cell_6t
Xbit_r90_c69 bl_69 br_69 wl_90 vdd gnd cell_6t
Xbit_r91_c69 bl_69 br_69 wl_91 vdd gnd cell_6t
Xbit_r92_c69 bl_69 br_69 wl_92 vdd gnd cell_6t
Xbit_r93_c69 bl_69 br_69 wl_93 vdd gnd cell_6t
Xbit_r94_c69 bl_69 br_69 wl_94 vdd gnd cell_6t
Xbit_r95_c69 bl_69 br_69 wl_95 vdd gnd cell_6t
Xbit_r96_c69 bl_69 br_69 wl_96 vdd gnd cell_6t
Xbit_r97_c69 bl_69 br_69 wl_97 vdd gnd cell_6t
Xbit_r98_c69 bl_69 br_69 wl_98 vdd gnd cell_6t
Xbit_r99_c69 bl_69 br_69 wl_99 vdd gnd cell_6t
Xbit_r100_c69 bl_69 br_69 wl_100 vdd gnd cell_6t
Xbit_r101_c69 bl_69 br_69 wl_101 vdd gnd cell_6t
Xbit_r102_c69 bl_69 br_69 wl_102 vdd gnd cell_6t
Xbit_r103_c69 bl_69 br_69 wl_103 vdd gnd cell_6t
Xbit_r104_c69 bl_69 br_69 wl_104 vdd gnd cell_6t
Xbit_r105_c69 bl_69 br_69 wl_105 vdd gnd cell_6t
Xbit_r106_c69 bl_69 br_69 wl_106 vdd gnd cell_6t
Xbit_r107_c69 bl_69 br_69 wl_107 vdd gnd cell_6t
Xbit_r108_c69 bl_69 br_69 wl_108 vdd gnd cell_6t
Xbit_r109_c69 bl_69 br_69 wl_109 vdd gnd cell_6t
Xbit_r110_c69 bl_69 br_69 wl_110 vdd gnd cell_6t
Xbit_r111_c69 bl_69 br_69 wl_111 vdd gnd cell_6t
Xbit_r112_c69 bl_69 br_69 wl_112 vdd gnd cell_6t
Xbit_r113_c69 bl_69 br_69 wl_113 vdd gnd cell_6t
Xbit_r114_c69 bl_69 br_69 wl_114 vdd gnd cell_6t
Xbit_r115_c69 bl_69 br_69 wl_115 vdd gnd cell_6t
Xbit_r116_c69 bl_69 br_69 wl_116 vdd gnd cell_6t
Xbit_r117_c69 bl_69 br_69 wl_117 vdd gnd cell_6t
Xbit_r118_c69 bl_69 br_69 wl_118 vdd gnd cell_6t
Xbit_r119_c69 bl_69 br_69 wl_119 vdd gnd cell_6t
Xbit_r120_c69 bl_69 br_69 wl_120 vdd gnd cell_6t
Xbit_r121_c69 bl_69 br_69 wl_121 vdd gnd cell_6t
Xbit_r122_c69 bl_69 br_69 wl_122 vdd gnd cell_6t
Xbit_r123_c69 bl_69 br_69 wl_123 vdd gnd cell_6t
Xbit_r124_c69 bl_69 br_69 wl_124 vdd gnd cell_6t
Xbit_r125_c69 bl_69 br_69 wl_125 vdd gnd cell_6t
Xbit_r126_c69 bl_69 br_69 wl_126 vdd gnd cell_6t
Xbit_r127_c69 bl_69 br_69 wl_127 vdd gnd cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd cell_6t
Xbit_r1_c70 bl_70 br_70 wl_1 vdd gnd cell_6t
Xbit_r2_c70 bl_70 br_70 wl_2 vdd gnd cell_6t
Xbit_r3_c70 bl_70 br_70 wl_3 vdd gnd cell_6t
Xbit_r4_c70 bl_70 br_70 wl_4 vdd gnd cell_6t
Xbit_r5_c70 bl_70 br_70 wl_5 vdd gnd cell_6t
Xbit_r6_c70 bl_70 br_70 wl_6 vdd gnd cell_6t
Xbit_r7_c70 bl_70 br_70 wl_7 vdd gnd cell_6t
Xbit_r8_c70 bl_70 br_70 wl_8 vdd gnd cell_6t
Xbit_r9_c70 bl_70 br_70 wl_9 vdd gnd cell_6t
Xbit_r10_c70 bl_70 br_70 wl_10 vdd gnd cell_6t
Xbit_r11_c70 bl_70 br_70 wl_11 vdd gnd cell_6t
Xbit_r12_c70 bl_70 br_70 wl_12 vdd gnd cell_6t
Xbit_r13_c70 bl_70 br_70 wl_13 vdd gnd cell_6t
Xbit_r14_c70 bl_70 br_70 wl_14 vdd gnd cell_6t
Xbit_r15_c70 bl_70 br_70 wl_15 vdd gnd cell_6t
Xbit_r16_c70 bl_70 br_70 wl_16 vdd gnd cell_6t
Xbit_r17_c70 bl_70 br_70 wl_17 vdd gnd cell_6t
Xbit_r18_c70 bl_70 br_70 wl_18 vdd gnd cell_6t
Xbit_r19_c70 bl_70 br_70 wl_19 vdd gnd cell_6t
Xbit_r20_c70 bl_70 br_70 wl_20 vdd gnd cell_6t
Xbit_r21_c70 bl_70 br_70 wl_21 vdd gnd cell_6t
Xbit_r22_c70 bl_70 br_70 wl_22 vdd gnd cell_6t
Xbit_r23_c70 bl_70 br_70 wl_23 vdd gnd cell_6t
Xbit_r24_c70 bl_70 br_70 wl_24 vdd gnd cell_6t
Xbit_r25_c70 bl_70 br_70 wl_25 vdd gnd cell_6t
Xbit_r26_c70 bl_70 br_70 wl_26 vdd gnd cell_6t
Xbit_r27_c70 bl_70 br_70 wl_27 vdd gnd cell_6t
Xbit_r28_c70 bl_70 br_70 wl_28 vdd gnd cell_6t
Xbit_r29_c70 bl_70 br_70 wl_29 vdd gnd cell_6t
Xbit_r30_c70 bl_70 br_70 wl_30 vdd gnd cell_6t
Xbit_r31_c70 bl_70 br_70 wl_31 vdd gnd cell_6t
Xbit_r32_c70 bl_70 br_70 wl_32 vdd gnd cell_6t
Xbit_r33_c70 bl_70 br_70 wl_33 vdd gnd cell_6t
Xbit_r34_c70 bl_70 br_70 wl_34 vdd gnd cell_6t
Xbit_r35_c70 bl_70 br_70 wl_35 vdd gnd cell_6t
Xbit_r36_c70 bl_70 br_70 wl_36 vdd gnd cell_6t
Xbit_r37_c70 bl_70 br_70 wl_37 vdd gnd cell_6t
Xbit_r38_c70 bl_70 br_70 wl_38 vdd gnd cell_6t
Xbit_r39_c70 bl_70 br_70 wl_39 vdd gnd cell_6t
Xbit_r40_c70 bl_70 br_70 wl_40 vdd gnd cell_6t
Xbit_r41_c70 bl_70 br_70 wl_41 vdd gnd cell_6t
Xbit_r42_c70 bl_70 br_70 wl_42 vdd gnd cell_6t
Xbit_r43_c70 bl_70 br_70 wl_43 vdd gnd cell_6t
Xbit_r44_c70 bl_70 br_70 wl_44 vdd gnd cell_6t
Xbit_r45_c70 bl_70 br_70 wl_45 vdd gnd cell_6t
Xbit_r46_c70 bl_70 br_70 wl_46 vdd gnd cell_6t
Xbit_r47_c70 bl_70 br_70 wl_47 vdd gnd cell_6t
Xbit_r48_c70 bl_70 br_70 wl_48 vdd gnd cell_6t
Xbit_r49_c70 bl_70 br_70 wl_49 vdd gnd cell_6t
Xbit_r50_c70 bl_70 br_70 wl_50 vdd gnd cell_6t
Xbit_r51_c70 bl_70 br_70 wl_51 vdd gnd cell_6t
Xbit_r52_c70 bl_70 br_70 wl_52 vdd gnd cell_6t
Xbit_r53_c70 bl_70 br_70 wl_53 vdd gnd cell_6t
Xbit_r54_c70 bl_70 br_70 wl_54 vdd gnd cell_6t
Xbit_r55_c70 bl_70 br_70 wl_55 vdd gnd cell_6t
Xbit_r56_c70 bl_70 br_70 wl_56 vdd gnd cell_6t
Xbit_r57_c70 bl_70 br_70 wl_57 vdd gnd cell_6t
Xbit_r58_c70 bl_70 br_70 wl_58 vdd gnd cell_6t
Xbit_r59_c70 bl_70 br_70 wl_59 vdd gnd cell_6t
Xbit_r60_c70 bl_70 br_70 wl_60 vdd gnd cell_6t
Xbit_r61_c70 bl_70 br_70 wl_61 vdd gnd cell_6t
Xbit_r62_c70 bl_70 br_70 wl_62 vdd gnd cell_6t
Xbit_r63_c70 bl_70 br_70 wl_63 vdd gnd cell_6t
Xbit_r64_c70 bl_70 br_70 wl_64 vdd gnd cell_6t
Xbit_r65_c70 bl_70 br_70 wl_65 vdd gnd cell_6t
Xbit_r66_c70 bl_70 br_70 wl_66 vdd gnd cell_6t
Xbit_r67_c70 bl_70 br_70 wl_67 vdd gnd cell_6t
Xbit_r68_c70 bl_70 br_70 wl_68 vdd gnd cell_6t
Xbit_r69_c70 bl_70 br_70 wl_69 vdd gnd cell_6t
Xbit_r70_c70 bl_70 br_70 wl_70 vdd gnd cell_6t
Xbit_r71_c70 bl_70 br_70 wl_71 vdd gnd cell_6t
Xbit_r72_c70 bl_70 br_70 wl_72 vdd gnd cell_6t
Xbit_r73_c70 bl_70 br_70 wl_73 vdd gnd cell_6t
Xbit_r74_c70 bl_70 br_70 wl_74 vdd gnd cell_6t
Xbit_r75_c70 bl_70 br_70 wl_75 vdd gnd cell_6t
Xbit_r76_c70 bl_70 br_70 wl_76 vdd gnd cell_6t
Xbit_r77_c70 bl_70 br_70 wl_77 vdd gnd cell_6t
Xbit_r78_c70 bl_70 br_70 wl_78 vdd gnd cell_6t
Xbit_r79_c70 bl_70 br_70 wl_79 vdd gnd cell_6t
Xbit_r80_c70 bl_70 br_70 wl_80 vdd gnd cell_6t
Xbit_r81_c70 bl_70 br_70 wl_81 vdd gnd cell_6t
Xbit_r82_c70 bl_70 br_70 wl_82 vdd gnd cell_6t
Xbit_r83_c70 bl_70 br_70 wl_83 vdd gnd cell_6t
Xbit_r84_c70 bl_70 br_70 wl_84 vdd gnd cell_6t
Xbit_r85_c70 bl_70 br_70 wl_85 vdd gnd cell_6t
Xbit_r86_c70 bl_70 br_70 wl_86 vdd gnd cell_6t
Xbit_r87_c70 bl_70 br_70 wl_87 vdd gnd cell_6t
Xbit_r88_c70 bl_70 br_70 wl_88 vdd gnd cell_6t
Xbit_r89_c70 bl_70 br_70 wl_89 vdd gnd cell_6t
Xbit_r90_c70 bl_70 br_70 wl_90 vdd gnd cell_6t
Xbit_r91_c70 bl_70 br_70 wl_91 vdd gnd cell_6t
Xbit_r92_c70 bl_70 br_70 wl_92 vdd gnd cell_6t
Xbit_r93_c70 bl_70 br_70 wl_93 vdd gnd cell_6t
Xbit_r94_c70 bl_70 br_70 wl_94 vdd gnd cell_6t
Xbit_r95_c70 bl_70 br_70 wl_95 vdd gnd cell_6t
Xbit_r96_c70 bl_70 br_70 wl_96 vdd gnd cell_6t
Xbit_r97_c70 bl_70 br_70 wl_97 vdd gnd cell_6t
Xbit_r98_c70 bl_70 br_70 wl_98 vdd gnd cell_6t
Xbit_r99_c70 bl_70 br_70 wl_99 vdd gnd cell_6t
Xbit_r100_c70 bl_70 br_70 wl_100 vdd gnd cell_6t
Xbit_r101_c70 bl_70 br_70 wl_101 vdd gnd cell_6t
Xbit_r102_c70 bl_70 br_70 wl_102 vdd gnd cell_6t
Xbit_r103_c70 bl_70 br_70 wl_103 vdd gnd cell_6t
Xbit_r104_c70 bl_70 br_70 wl_104 vdd gnd cell_6t
Xbit_r105_c70 bl_70 br_70 wl_105 vdd gnd cell_6t
Xbit_r106_c70 bl_70 br_70 wl_106 vdd gnd cell_6t
Xbit_r107_c70 bl_70 br_70 wl_107 vdd gnd cell_6t
Xbit_r108_c70 bl_70 br_70 wl_108 vdd gnd cell_6t
Xbit_r109_c70 bl_70 br_70 wl_109 vdd gnd cell_6t
Xbit_r110_c70 bl_70 br_70 wl_110 vdd gnd cell_6t
Xbit_r111_c70 bl_70 br_70 wl_111 vdd gnd cell_6t
Xbit_r112_c70 bl_70 br_70 wl_112 vdd gnd cell_6t
Xbit_r113_c70 bl_70 br_70 wl_113 vdd gnd cell_6t
Xbit_r114_c70 bl_70 br_70 wl_114 vdd gnd cell_6t
Xbit_r115_c70 bl_70 br_70 wl_115 vdd gnd cell_6t
Xbit_r116_c70 bl_70 br_70 wl_116 vdd gnd cell_6t
Xbit_r117_c70 bl_70 br_70 wl_117 vdd gnd cell_6t
Xbit_r118_c70 bl_70 br_70 wl_118 vdd gnd cell_6t
Xbit_r119_c70 bl_70 br_70 wl_119 vdd gnd cell_6t
Xbit_r120_c70 bl_70 br_70 wl_120 vdd gnd cell_6t
Xbit_r121_c70 bl_70 br_70 wl_121 vdd gnd cell_6t
Xbit_r122_c70 bl_70 br_70 wl_122 vdd gnd cell_6t
Xbit_r123_c70 bl_70 br_70 wl_123 vdd gnd cell_6t
Xbit_r124_c70 bl_70 br_70 wl_124 vdd gnd cell_6t
Xbit_r125_c70 bl_70 br_70 wl_125 vdd gnd cell_6t
Xbit_r126_c70 bl_70 br_70 wl_126 vdd gnd cell_6t
Xbit_r127_c70 bl_70 br_70 wl_127 vdd gnd cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd cell_6t
Xbit_r1_c71 bl_71 br_71 wl_1 vdd gnd cell_6t
Xbit_r2_c71 bl_71 br_71 wl_2 vdd gnd cell_6t
Xbit_r3_c71 bl_71 br_71 wl_3 vdd gnd cell_6t
Xbit_r4_c71 bl_71 br_71 wl_4 vdd gnd cell_6t
Xbit_r5_c71 bl_71 br_71 wl_5 vdd gnd cell_6t
Xbit_r6_c71 bl_71 br_71 wl_6 vdd gnd cell_6t
Xbit_r7_c71 bl_71 br_71 wl_7 vdd gnd cell_6t
Xbit_r8_c71 bl_71 br_71 wl_8 vdd gnd cell_6t
Xbit_r9_c71 bl_71 br_71 wl_9 vdd gnd cell_6t
Xbit_r10_c71 bl_71 br_71 wl_10 vdd gnd cell_6t
Xbit_r11_c71 bl_71 br_71 wl_11 vdd gnd cell_6t
Xbit_r12_c71 bl_71 br_71 wl_12 vdd gnd cell_6t
Xbit_r13_c71 bl_71 br_71 wl_13 vdd gnd cell_6t
Xbit_r14_c71 bl_71 br_71 wl_14 vdd gnd cell_6t
Xbit_r15_c71 bl_71 br_71 wl_15 vdd gnd cell_6t
Xbit_r16_c71 bl_71 br_71 wl_16 vdd gnd cell_6t
Xbit_r17_c71 bl_71 br_71 wl_17 vdd gnd cell_6t
Xbit_r18_c71 bl_71 br_71 wl_18 vdd gnd cell_6t
Xbit_r19_c71 bl_71 br_71 wl_19 vdd gnd cell_6t
Xbit_r20_c71 bl_71 br_71 wl_20 vdd gnd cell_6t
Xbit_r21_c71 bl_71 br_71 wl_21 vdd gnd cell_6t
Xbit_r22_c71 bl_71 br_71 wl_22 vdd gnd cell_6t
Xbit_r23_c71 bl_71 br_71 wl_23 vdd gnd cell_6t
Xbit_r24_c71 bl_71 br_71 wl_24 vdd gnd cell_6t
Xbit_r25_c71 bl_71 br_71 wl_25 vdd gnd cell_6t
Xbit_r26_c71 bl_71 br_71 wl_26 vdd gnd cell_6t
Xbit_r27_c71 bl_71 br_71 wl_27 vdd gnd cell_6t
Xbit_r28_c71 bl_71 br_71 wl_28 vdd gnd cell_6t
Xbit_r29_c71 bl_71 br_71 wl_29 vdd gnd cell_6t
Xbit_r30_c71 bl_71 br_71 wl_30 vdd gnd cell_6t
Xbit_r31_c71 bl_71 br_71 wl_31 vdd gnd cell_6t
Xbit_r32_c71 bl_71 br_71 wl_32 vdd gnd cell_6t
Xbit_r33_c71 bl_71 br_71 wl_33 vdd gnd cell_6t
Xbit_r34_c71 bl_71 br_71 wl_34 vdd gnd cell_6t
Xbit_r35_c71 bl_71 br_71 wl_35 vdd gnd cell_6t
Xbit_r36_c71 bl_71 br_71 wl_36 vdd gnd cell_6t
Xbit_r37_c71 bl_71 br_71 wl_37 vdd gnd cell_6t
Xbit_r38_c71 bl_71 br_71 wl_38 vdd gnd cell_6t
Xbit_r39_c71 bl_71 br_71 wl_39 vdd gnd cell_6t
Xbit_r40_c71 bl_71 br_71 wl_40 vdd gnd cell_6t
Xbit_r41_c71 bl_71 br_71 wl_41 vdd gnd cell_6t
Xbit_r42_c71 bl_71 br_71 wl_42 vdd gnd cell_6t
Xbit_r43_c71 bl_71 br_71 wl_43 vdd gnd cell_6t
Xbit_r44_c71 bl_71 br_71 wl_44 vdd gnd cell_6t
Xbit_r45_c71 bl_71 br_71 wl_45 vdd gnd cell_6t
Xbit_r46_c71 bl_71 br_71 wl_46 vdd gnd cell_6t
Xbit_r47_c71 bl_71 br_71 wl_47 vdd gnd cell_6t
Xbit_r48_c71 bl_71 br_71 wl_48 vdd gnd cell_6t
Xbit_r49_c71 bl_71 br_71 wl_49 vdd gnd cell_6t
Xbit_r50_c71 bl_71 br_71 wl_50 vdd gnd cell_6t
Xbit_r51_c71 bl_71 br_71 wl_51 vdd gnd cell_6t
Xbit_r52_c71 bl_71 br_71 wl_52 vdd gnd cell_6t
Xbit_r53_c71 bl_71 br_71 wl_53 vdd gnd cell_6t
Xbit_r54_c71 bl_71 br_71 wl_54 vdd gnd cell_6t
Xbit_r55_c71 bl_71 br_71 wl_55 vdd gnd cell_6t
Xbit_r56_c71 bl_71 br_71 wl_56 vdd gnd cell_6t
Xbit_r57_c71 bl_71 br_71 wl_57 vdd gnd cell_6t
Xbit_r58_c71 bl_71 br_71 wl_58 vdd gnd cell_6t
Xbit_r59_c71 bl_71 br_71 wl_59 vdd gnd cell_6t
Xbit_r60_c71 bl_71 br_71 wl_60 vdd gnd cell_6t
Xbit_r61_c71 bl_71 br_71 wl_61 vdd gnd cell_6t
Xbit_r62_c71 bl_71 br_71 wl_62 vdd gnd cell_6t
Xbit_r63_c71 bl_71 br_71 wl_63 vdd gnd cell_6t
Xbit_r64_c71 bl_71 br_71 wl_64 vdd gnd cell_6t
Xbit_r65_c71 bl_71 br_71 wl_65 vdd gnd cell_6t
Xbit_r66_c71 bl_71 br_71 wl_66 vdd gnd cell_6t
Xbit_r67_c71 bl_71 br_71 wl_67 vdd gnd cell_6t
Xbit_r68_c71 bl_71 br_71 wl_68 vdd gnd cell_6t
Xbit_r69_c71 bl_71 br_71 wl_69 vdd gnd cell_6t
Xbit_r70_c71 bl_71 br_71 wl_70 vdd gnd cell_6t
Xbit_r71_c71 bl_71 br_71 wl_71 vdd gnd cell_6t
Xbit_r72_c71 bl_71 br_71 wl_72 vdd gnd cell_6t
Xbit_r73_c71 bl_71 br_71 wl_73 vdd gnd cell_6t
Xbit_r74_c71 bl_71 br_71 wl_74 vdd gnd cell_6t
Xbit_r75_c71 bl_71 br_71 wl_75 vdd gnd cell_6t
Xbit_r76_c71 bl_71 br_71 wl_76 vdd gnd cell_6t
Xbit_r77_c71 bl_71 br_71 wl_77 vdd gnd cell_6t
Xbit_r78_c71 bl_71 br_71 wl_78 vdd gnd cell_6t
Xbit_r79_c71 bl_71 br_71 wl_79 vdd gnd cell_6t
Xbit_r80_c71 bl_71 br_71 wl_80 vdd gnd cell_6t
Xbit_r81_c71 bl_71 br_71 wl_81 vdd gnd cell_6t
Xbit_r82_c71 bl_71 br_71 wl_82 vdd gnd cell_6t
Xbit_r83_c71 bl_71 br_71 wl_83 vdd gnd cell_6t
Xbit_r84_c71 bl_71 br_71 wl_84 vdd gnd cell_6t
Xbit_r85_c71 bl_71 br_71 wl_85 vdd gnd cell_6t
Xbit_r86_c71 bl_71 br_71 wl_86 vdd gnd cell_6t
Xbit_r87_c71 bl_71 br_71 wl_87 vdd gnd cell_6t
Xbit_r88_c71 bl_71 br_71 wl_88 vdd gnd cell_6t
Xbit_r89_c71 bl_71 br_71 wl_89 vdd gnd cell_6t
Xbit_r90_c71 bl_71 br_71 wl_90 vdd gnd cell_6t
Xbit_r91_c71 bl_71 br_71 wl_91 vdd gnd cell_6t
Xbit_r92_c71 bl_71 br_71 wl_92 vdd gnd cell_6t
Xbit_r93_c71 bl_71 br_71 wl_93 vdd gnd cell_6t
Xbit_r94_c71 bl_71 br_71 wl_94 vdd gnd cell_6t
Xbit_r95_c71 bl_71 br_71 wl_95 vdd gnd cell_6t
Xbit_r96_c71 bl_71 br_71 wl_96 vdd gnd cell_6t
Xbit_r97_c71 bl_71 br_71 wl_97 vdd gnd cell_6t
Xbit_r98_c71 bl_71 br_71 wl_98 vdd gnd cell_6t
Xbit_r99_c71 bl_71 br_71 wl_99 vdd gnd cell_6t
Xbit_r100_c71 bl_71 br_71 wl_100 vdd gnd cell_6t
Xbit_r101_c71 bl_71 br_71 wl_101 vdd gnd cell_6t
Xbit_r102_c71 bl_71 br_71 wl_102 vdd gnd cell_6t
Xbit_r103_c71 bl_71 br_71 wl_103 vdd gnd cell_6t
Xbit_r104_c71 bl_71 br_71 wl_104 vdd gnd cell_6t
Xbit_r105_c71 bl_71 br_71 wl_105 vdd gnd cell_6t
Xbit_r106_c71 bl_71 br_71 wl_106 vdd gnd cell_6t
Xbit_r107_c71 bl_71 br_71 wl_107 vdd gnd cell_6t
Xbit_r108_c71 bl_71 br_71 wl_108 vdd gnd cell_6t
Xbit_r109_c71 bl_71 br_71 wl_109 vdd gnd cell_6t
Xbit_r110_c71 bl_71 br_71 wl_110 vdd gnd cell_6t
Xbit_r111_c71 bl_71 br_71 wl_111 vdd gnd cell_6t
Xbit_r112_c71 bl_71 br_71 wl_112 vdd gnd cell_6t
Xbit_r113_c71 bl_71 br_71 wl_113 vdd gnd cell_6t
Xbit_r114_c71 bl_71 br_71 wl_114 vdd gnd cell_6t
Xbit_r115_c71 bl_71 br_71 wl_115 vdd gnd cell_6t
Xbit_r116_c71 bl_71 br_71 wl_116 vdd gnd cell_6t
Xbit_r117_c71 bl_71 br_71 wl_117 vdd gnd cell_6t
Xbit_r118_c71 bl_71 br_71 wl_118 vdd gnd cell_6t
Xbit_r119_c71 bl_71 br_71 wl_119 vdd gnd cell_6t
Xbit_r120_c71 bl_71 br_71 wl_120 vdd gnd cell_6t
Xbit_r121_c71 bl_71 br_71 wl_121 vdd gnd cell_6t
Xbit_r122_c71 bl_71 br_71 wl_122 vdd gnd cell_6t
Xbit_r123_c71 bl_71 br_71 wl_123 vdd gnd cell_6t
Xbit_r124_c71 bl_71 br_71 wl_124 vdd gnd cell_6t
Xbit_r125_c71 bl_71 br_71 wl_125 vdd gnd cell_6t
Xbit_r126_c71 bl_71 br_71 wl_126 vdd gnd cell_6t
Xbit_r127_c71 bl_71 br_71 wl_127 vdd gnd cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd cell_6t
Xbit_r1_c72 bl_72 br_72 wl_1 vdd gnd cell_6t
Xbit_r2_c72 bl_72 br_72 wl_2 vdd gnd cell_6t
Xbit_r3_c72 bl_72 br_72 wl_3 vdd gnd cell_6t
Xbit_r4_c72 bl_72 br_72 wl_4 vdd gnd cell_6t
Xbit_r5_c72 bl_72 br_72 wl_5 vdd gnd cell_6t
Xbit_r6_c72 bl_72 br_72 wl_6 vdd gnd cell_6t
Xbit_r7_c72 bl_72 br_72 wl_7 vdd gnd cell_6t
Xbit_r8_c72 bl_72 br_72 wl_8 vdd gnd cell_6t
Xbit_r9_c72 bl_72 br_72 wl_9 vdd gnd cell_6t
Xbit_r10_c72 bl_72 br_72 wl_10 vdd gnd cell_6t
Xbit_r11_c72 bl_72 br_72 wl_11 vdd gnd cell_6t
Xbit_r12_c72 bl_72 br_72 wl_12 vdd gnd cell_6t
Xbit_r13_c72 bl_72 br_72 wl_13 vdd gnd cell_6t
Xbit_r14_c72 bl_72 br_72 wl_14 vdd gnd cell_6t
Xbit_r15_c72 bl_72 br_72 wl_15 vdd gnd cell_6t
Xbit_r16_c72 bl_72 br_72 wl_16 vdd gnd cell_6t
Xbit_r17_c72 bl_72 br_72 wl_17 vdd gnd cell_6t
Xbit_r18_c72 bl_72 br_72 wl_18 vdd gnd cell_6t
Xbit_r19_c72 bl_72 br_72 wl_19 vdd gnd cell_6t
Xbit_r20_c72 bl_72 br_72 wl_20 vdd gnd cell_6t
Xbit_r21_c72 bl_72 br_72 wl_21 vdd gnd cell_6t
Xbit_r22_c72 bl_72 br_72 wl_22 vdd gnd cell_6t
Xbit_r23_c72 bl_72 br_72 wl_23 vdd gnd cell_6t
Xbit_r24_c72 bl_72 br_72 wl_24 vdd gnd cell_6t
Xbit_r25_c72 bl_72 br_72 wl_25 vdd gnd cell_6t
Xbit_r26_c72 bl_72 br_72 wl_26 vdd gnd cell_6t
Xbit_r27_c72 bl_72 br_72 wl_27 vdd gnd cell_6t
Xbit_r28_c72 bl_72 br_72 wl_28 vdd gnd cell_6t
Xbit_r29_c72 bl_72 br_72 wl_29 vdd gnd cell_6t
Xbit_r30_c72 bl_72 br_72 wl_30 vdd gnd cell_6t
Xbit_r31_c72 bl_72 br_72 wl_31 vdd gnd cell_6t
Xbit_r32_c72 bl_72 br_72 wl_32 vdd gnd cell_6t
Xbit_r33_c72 bl_72 br_72 wl_33 vdd gnd cell_6t
Xbit_r34_c72 bl_72 br_72 wl_34 vdd gnd cell_6t
Xbit_r35_c72 bl_72 br_72 wl_35 vdd gnd cell_6t
Xbit_r36_c72 bl_72 br_72 wl_36 vdd gnd cell_6t
Xbit_r37_c72 bl_72 br_72 wl_37 vdd gnd cell_6t
Xbit_r38_c72 bl_72 br_72 wl_38 vdd gnd cell_6t
Xbit_r39_c72 bl_72 br_72 wl_39 vdd gnd cell_6t
Xbit_r40_c72 bl_72 br_72 wl_40 vdd gnd cell_6t
Xbit_r41_c72 bl_72 br_72 wl_41 vdd gnd cell_6t
Xbit_r42_c72 bl_72 br_72 wl_42 vdd gnd cell_6t
Xbit_r43_c72 bl_72 br_72 wl_43 vdd gnd cell_6t
Xbit_r44_c72 bl_72 br_72 wl_44 vdd gnd cell_6t
Xbit_r45_c72 bl_72 br_72 wl_45 vdd gnd cell_6t
Xbit_r46_c72 bl_72 br_72 wl_46 vdd gnd cell_6t
Xbit_r47_c72 bl_72 br_72 wl_47 vdd gnd cell_6t
Xbit_r48_c72 bl_72 br_72 wl_48 vdd gnd cell_6t
Xbit_r49_c72 bl_72 br_72 wl_49 vdd gnd cell_6t
Xbit_r50_c72 bl_72 br_72 wl_50 vdd gnd cell_6t
Xbit_r51_c72 bl_72 br_72 wl_51 vdd gnd cell_6t
Xbit_r52_c72 bl_72 br_72 wl_52 vdd gnd cell_6t
Xbit_r53_c72 bl_72 br_72 wl_53 vdd gnd cell_6t
Xbit_r54_c72 bl_72 br_72 wl_54 vdd gnd cell_6t
Xbit_r55_c72 bl_72 br_72 wl_55 vdd gnd cell_6t
Xbit_r56_c72 bl_72 br_72 wl_56 vdd gnd cell_6t
Xbit_r57_c72 bl_72 br_72 wl_57 vdd gnd cell_6t
Xbit_r58_c72 bl_72 br_72 wl_58 vdd gnd cell_6t
Xbit_r59_c72 bl_72 br_72 wl_59 vdd gnd cell_6t
Xbit_r60_c72 bl_72 br_72 wl_60 vdd gnd cell_6t
Xbit_r61_c72 bl_72 br_72 wl_61 vdd gnd cell_6t
Xbit_r62_c72 bl_72 br_72 wl_62 vdd gnd cell_6t
Xbit_r63_c72 bl_72 br_72 wl_63 vdd gnd cell_6t
Xbit_r64_c72 bl_72 br_72 wl_64 vdd gnd cell_6t
Xbit_r65_c72 bl_72 br_72 wl_65 vdd gnd cell_6t
Xbit_r66_c72 bl_72 br_72 wl_66 vdd gnd cell_6t
Xbit_r67_c72 bl_72 br_72 wl_67 vdd gnd cell_6t
Xbit_r68_c72 bl_72 br_72 wl_68 vdd gnd cell_6t
Xbit_r69_c72 bl_72 br_72 wl_69 vdd gnd cell_6t
Xbit_r70_c72 bl_72 br_72 wl_70 vdd gnd cell_6t
Xbit_r71_c72 bl_72 br_72 wl_71 vdd gnd cell_6t
Xbit_r72_c72 bl_72 br_72 wl_72 vdd gnd cell_6t
Xbit_r73_c72 bl_72 br_72 wl_73 vdd gnd cell_6t
Xbit_r74_c72 bl_72 br_72 wl_74 vdd gnd cell_6t
Xbit_r75_c72 bl_72 br_72 wl_75 vdd gnd cell_6t
Xbit_r76_c72 bl_72 br_72 wl_76 vdd gnd cell_6t
Xbit_r77_c72 bl_72 br_72 wl_77 vdd gnd cell_6t
Xbit_r78_c72 bl_72 br_72 wl_78 vdd gnd cell_6t
Xbit_r79_c72 bl_72 br_72 wl_79 vdd gnd cell_6t
Xbit_r80_c72 bl_72 br_72 wl_80 vdd gnd cell_6t
Xbit_r81_c72 bl_72 br_72 wl_81 vdd gnd cell_6t
Xbit_r82_c72 bl_72 br_72 wl_82 vdd gnd cell_6t
Xbit_r83_c72 bl_72 br_72 wl_83 vdd gnd cell_6t
Xbit_r84_c72 bl_72 br_72 wl_84 vdd gnd cell_6t
Xbit_r85_c72 bl_72 br_72 wl_85 vdd gnd cell_6t
Xbit_r86_c72 bl_72 br_72 wl_86 vdd gnd cell_6t
Xbit_r87_c72 bl_72 br_72 wl_87 vdd gnd cell_6t
Xbit_r88_c72 bl_72 br_72 wl_88 vdd gnd cell_6t
Xbit_r89_c72 bl_72 br_72 wl_89 vdd gnd cell_6t
Xbit_r90_c72 bl_72 br_72 wl_90 vdd gnd cell_6t
Xbit_r91_c72 bl_72 br_72 wl_91 vdd gnd cell_6t
Xbit_r92_c72 bl_72 br_72 wl_92 vdd gnd cell_6t
Xbit_r93_c72 bl_72 br_72 wl_93 vdd gnd cell_6t
Xbit_r94_c72 bl_72 br_72 wl_94 vdd gnd cell_6t
Xbit_r95_c72 bl_72 br_72 wl_95 vdd gnd cell_6t
Xbit_r96_c72 bl_72 br_72 wl_96 vdd gnd cell_6t
Xbit_r97_c72 bl_72 br_72 wl_97 vdd gnd cell_6t
Xbit_r98_c72 bl_72 br_72 wl_98 vdd gnd cell_6t
Xbit_r99_c72 bl_72 br_72 wl_99 vdd gnd cell_6t
Xbit_r100_c72 bl_72 br_72 wl_100 vdd gnd cell_6t
Xbit_r101_c72 bl_72 br_72 wl_101 vdd gnd cell_6t
Xbit_r102_c72 bl_72 br_72 wl_102 vdd gnd cell_6t
Xbit_r103_c72 bl_72 br_72 wl_103 vdd gnd cell_6t
Xbit_r104_c72 bl_72 br_72 wl_104 vdd gnd cell_6t
Xbit_r105_c72 bl_72 br_72 wl_105 vdd gnd cell_6t
Xbit_r106_c72 bl_72 br_72 wl_106 vdd gnd cell_6t
Xbit_r107_c72 bl_72 br_72 wl_107 vdd gnd cell_6t
Xbit_r108_c72 bl_72 br_72 wl_108 vdd gnd cell_6t
Xbit_r109_c72 bl_72 br_72 wl_109 vdd gnd cell_6t
Xbit_r110_c72 bl_72 br_72 wl_110 vdd gnd cell_6t
Xbit_r111_c72 bl_72 br_72 wl_111 vdd gnd cell_6t
Xbit_r112_c72 bl_72 br_72 wl_112 vdd gnd cell_6t
Xbit_r113_c72 bl_72 br_72 wl_113 vdd gnd cell_6t
Xbit_r114_c72 bl_72 br_72 wl_114 vdd gnd cell_6t
Xbit_r115_c72 bl_72 br_72 wl_115 vdd gnd cell_6t
Xbit_r116_c72 bl_72 br_72 wl_116 vdd gnd cell_6t
Xbit_r117_c72 bl_72 br_72 wl_117 vdd gnd cell_6t
Xbit_r118_c72 bl_72 br_72 wl_118 vdd gnd cell_6t
Xbit_r119_c72 bl_72 br_72 wl_119 vdd gnd cell_6t
Xbit_r120_c72 bl_72 br_72 wl_120 vdd gnd cell_6t
Xbit_r121_c72 bl_72 br_72 wl_121 vdd gnd cell_6t
Xbit_r122_c72 bl_72 br_72 wl_122 vdd gnd cell_6t
Xbit_r123_c72 bl_72 br_72 wl_123 vdd gnd cell_6t
Xbit_r124_c72 bl_72 br_72 wl_124 vdd gnd cell_6t
Xbit_r125_c72 bl_72 br_72 wl_125 vdd gnd cell_6t
Xbit_r126_c72 bl_72 br_72 wl_126 vdd gnd cell_6t
Xbit_r127_c72 bl_72 br_72 wl_127 vdd gnd cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd cell_6t
Xbit_r1_c73 bl_73 br_73 wl_1 vdd gnd cell_6t
Xbit_r2_c73 bl_73 br_73 wl_2 vdd gnd cell_6t
Xbit_r3_c73 bl_73 br_73 wl_3 vdd gnd cell_6t
Xbit_r4_c73 bl_73 br_73 wl_4 vdd gnd cell_6t
Xbit_r5_c73 bl_73 br_73 wl_5 vdd gnd cell_6t
Xbit_r6_c73 bl_73 br_73 wl_6 vdd gnd cell_6t
Xbit_r7_c73 bl_73 br_73 wl_7 vdd gnd cell_6t
Xbit_r8_c73 bl_73 br_73 wl_8 vdd gnd cell_6t
Xbit_r9_c73 bl_73 br_73 wl_9 vdd gnd cell_6t
Xbit_r10_c73 bl_73 br_73 wl_10 vdd gnd cell_6t
Xbit_r11_c73 bl_73 br_73 wl_11 vdd gnd cell_6t
Xbit_r12_c73 bl_73 br_73 wl_12 vdd gnd cell_6t
Xbit_r13_c73 bl_73 br_73 wl_13 vdd gnd cell_6t
Xbit_r14_c73 bl_73 br_73 wl_14 vdd gnd cell_6t
Xbit_r15_c73 bl_73 br_73 wl_15 vdd gnd cell_6t
Xbit_r16_c73 bl_73 br_73 wl_16 vdd gnd cell_6t
Xbit_r17_c73 bl_73 br_73 wl_17 vdd gnd cell_6t
Xbit_r18_c73 bl_73 br_73 wl_18 vdd gnd cell_6t
Xbit_r19_c73 bl_73 br_73 wl_19 vdd gnd cell_6t
Xbit_r20_c73 bl_73 br_73 wl_20 vdd gnd cell_6t
Xbit_r21_c73 bl_73 br_73 wl_21 vdd gnd cell_6t
Xbit_r22_c73 bl_73 br_73 wl_22 vdd gnd cell_6t
Xbit_r23_c73 bl_73 br_73 wl_23 vdd gnd cell_6t
Xbit_r24_c73 bl_73 br_73 wl_24 vdd gnd cell_6t
Xbit_r25_c73 bl_73 br_73 wl_25 vdd gnd cell_6t
Xbit_r26_c73 bl_73 br_73 wl_26 vdd gnd cell_6t
Xbit_r27_c73 bl_73 br_73 wl_27 vdd gnd cell_6t
Xbit_r28_c73 bl_73 br_73 wl_28 vdd gnd cell_6t
Xbit_r29_c73 bl_73 br_73 wl_29 vdd gnd cell_6t
Xbit_r30_c73 bl_73 br_73 wl_30 vdd gnd cell_6t
Xbit_r31_c73 bl_73 br_73 wl_31 vdd gnd cell_6t
Xbit_r32_c73 bl_73 br_73 wl_32 vdd gnd cell_6t
Xbit_r33_c73 bl_73 br_73 wl_33 vdd gnd cell_6t
Xbit_r34_c73 bl_73 br_73 wl_34 vdd gnd cell_6t
Xbit_r35_c73 bl_73 br_73 wl_35 vdd gnd cell_6t
Xbit_r36_c73 bl_73 br_73 wl_36 vdd gnd cell_6t
Xbit_r37_c73 bl_73 br_73 wl_37 vdd gnd cell_6t
Xbit_r38_c73 bl_73 br_73 wl_38 vdd gnd cell_6t
Xbit_r39_c73 bl_73 br_73 wl_39 vdd gnd cell_6t
Xbit_r40_c73 bl_73 br_73 wl_40 vdd gnd cell_6t
Xbit_r41_c73 bl_73 br_73 wl_41 vdd gnd cell_6t
Xbit_r42_c73 bl_73 br_73 wl_42 vdd gnd cell_6t
Xbit_r43_c73 bl_73 br_73 wl_43 vdd gnd cell_6t
Xbit_r44_c73 bl_73 br_73 wl_44 vdd gnd cell_6t
Xbit_r45_c73 bl_73 br_73 wl_45 vdd gnd cell_6t
Xbit_r46_c73 bl_73 br_73 wl_46 vdd gnd cell_6t
Xbit_r47_c73 bl_73 br_73 wl_47 vdd gnd cell_6t
Xbit_r48_c73 bl_73 br_73 wl_48 vdd gnd cell_6t
Xbit_r49_c73 bl_73 br_73 wl_49 vdd gnd cell_6t
Xbit_r50_c73 bl_73 br_73 wl_50 vdd gnd cell_6t
Xbit_r51_c73 bl_73 br_73 wl_51 vdd gnd cell_6t
Xbit_r52_c73 bl_73 br_73 wl_52 vdd gnd cell_6t
Xbit_r53_c73 bl_73 br_73 wl_53 vdd gnd cell_6t
Xbit_r54_c73 bl_73 br_73 wl_54 vdd gnd cell_6t
Xbit_r55_c73 bl_73 br_73 wl_55 vdd gnd cell_6t
Xbit_r56_c73 bl_73 br_73 wl_56 vdd gnd cell_6t
Xbit_r57_c73 bl_73 br_73 wl_57 vdd gnd cell_6t
Xbit_r58_c73 bl_73 br_73 wl_58 vdd gnd cell_6t
Xbit_r59_c73 bl_73 br_73 wl_59 vdd gnd cell_6t
Xbit_r60_c73 bl_73 br_73 wl_60 vdd gnd cell_6t
Xbit_r61_c73 bl_73 br_73 wl_61 vdd gnd cell_6t
Xbit_r62_c73 bl_73 br_73 wl_62 vdd gnd cell_6t
Xbit_r63_c73 bl_73 br_73 wl_63 vdd gnd cell_6t
Xbit_r64_c73 bl_73 br_73 wl_64 vdd gnd cell_6t
Xbit_r65_c73 bl_73 br_73 wl_65 vdd gnd cell_6t
Xbit_r66_c73 bl_73 br_73 wl_66 vdd gnd cell_6t
Xbit_r67_c73 bl_73 br_73 wl_67 vdd gnd cell_6t
Xbit_r68_c73 bl_73 br_73 wl_68 vdd gnd cell_6t
Xbit_r69_c73 bl_73 br_73 wl_69 vdd gnd cell_6t
Xbit_r70_c73 bl_73 br_73 wl_70 vdd gnd cell_6t
Xbit_r71_c73 bl_73 br_73 wl_71 vdd gnd cell_6t
Xbit_r72_c73 bl_73 br_73 wl_72 vdd gnd cell_6t
Xbit_r73_c73 bl_73 br_73 wl_73 vdd gnd cell_6t
Xbit_r74_c73 bl_73 br_73 wl_74 vdd gnd cell_6t
Xbit_r75_c73 bl_73 br_73 wl_75 vdd gnd cell_6t
Xbit_r76_c73 bl_73 br_73 wl_76 vdd gnd cell_6t
Xbit_r77_c73 bl_73 br_73 wl_77 vdd gnd cell_6t
Xbit_r78_c73 bl_73 br_73 wl_78 vdd gnd cell_6t
Xbit_r79_c73 bl_73 br_73 wl_79 vdd gnd cell_6t
Xbit_r80_c73 bl_73 br_73 wl_80 vdd gnd cell_6t
Xbit_r81_c73 bl_73 br_73 wl_81 vdd gnd cell_6t
Xbit_r82_c73 bl_73 br_73 wl_82 vdd gnd cell_6t
Xbit_r83_c73 bl_73 br_73 wl_83 vdd gnd cell_6t
Xbit_r84_c73 bl_73 br_73 wl_84 vdd gnd cell_6t
Xbit_r85_c73 bl_73 br_73 wl_85 vdd gnd cell_6t
Xbit_r86_c73 bl_73 br_73 wl_86 vdd gnd cell_6t
Xbit_r87_c73 bl_73 br_73 wl_87 vdd gnd cell_6t
Xbit_r88_c73 bl_73 br_73 wl_88 vdd gnd cell_6t
Xbit_r89_c73 bl_73 br_73 wl_89 vdd gnd cell_6t
Xbit_r90_c73 bl_73 br_73 wl_90 vdd gnd cell_6t
Xbit_r91_c73 bl_73 br_73 wl_91 vdd gnd cell_6t
Xbit_r92_c73 bl_73 br_73 wl_92 vdd gnd cell_6t
Xbit_r93_c73 bl_73 br_73 wl_93 vdd gnd cell_6t
Xbit_r94_c73 bl_73 br_73 wl_94 vdd gnd cell_6t
Xbit_r95_c73 bl_73 br_73 wl_95 vdd gnd cell_6t
Xbit_r96_c73 bl_73 br_73 wl_96 vdd gnd cell_6t
Xbit_r97_c73 bl_73 br_73 wl_97 vdd gnd cell_6t
Xbit_r98_c73 bl_73 br_73 wl_98 vdd gnd cell_6t
Xbit_r99_c73 bl_73 br_73 wl_99 vdd gnd cell_6t
Xbit_r100_c73 bl_73 br_73 wl_100 vdd gnd cell_6t
Xbit_r101_c73 bl_73 br_73 wl_101 vdd gnd cell_6t
Xbit_r102_c73 bl_73 br_73 wl_102 vdd gnd cell_6t
Xbit_r103_c73 bl_73 br_73 wl_103 vdd gnd cell_6t
Xbit_r104_c73 bl_73 br_73 wl_104 vdd gnd cell_6t
Xbit_r105_c73 bl_73 br_73 wl_105 vdd gnd cell_6t
Xbit_r106_c73 bl_73 br_73 wl_106 vdd gnd cell_6t
Xbit_r107_c73 bl_73 br_73 wl_107 vdd gnd cell_6t
Xbit_r108_c73 bl_73 br_73 wl_108 vdd gnd cell_6t
Xbit_r109_c73 bl_73 br_73 wl_109 vdd gnd cell_6t
Xbit_r110_c73 bl_73 br_73 wl_110 vdd gnd cell_6t
Xbit_r111_c73 bl_73 br_73 wl_111 vdd gnd cell_6t
Xbit_r112_c73 bl_73 br_73 wl_112 vdd gnd cell_6t
Xbit_r113_c73 bl_73 br_73 wl_113 vdd gnd cell_6t
Xbit_r114_c73 bl_73 br_73 wl_114 vdd gnd cell_6t
Xbit_r115_c73 bl_73 br_73 wl_115 vdd gnd cell_6t
Xbit_r116_c73 bl_73 br_73 wl_116 vdd gnd cell_6t
Xbit_r117_c73 bl_73 br_73 wl_117 vdd gnd cell_6t
Xbit_r118_c73 bl_73 br_73 wl_118 vdd gnd cell_6t
Xbit_r119_c73 bl_73 br_73 wl_119 vdd gnd cell_6t
Xbit_r120_c73 bl_73 br_73 wl_120 vdd gnd cell_6t
Xbit_r121_c73 bl_73 br_73 wl_121 vdd gnd cell_6t
Xbit_r122_c73 bl_73 br_73 wl_122 vdd gnd cell_6t
Xbit_r123_c73 bl_73 br_73 wl_123 vdd gnd cell_6t
Xbit_r124_c73 bl_73 br_73 wl_124 vdd gnd cell_6t
Xbit_r125_c73 bl_73 br_73 wl_125 vdd gnd cell_6t
Xbit_r126_c73 bl_73 br_73 wl_126 vdd gnd cell_6t
Xbit_r127_c73 bl_73 br_73 wl_127 vdd gnd cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd cell_6t
Xbit_r1_c74 bl_74 br_74 wl_1 vdd gnd cell_6t
Xbit_r2_c74 bl_74 br_74 wl_2 vdd gnd cell_6t
Xbit_r3_c74 bl_74 br_74 wl_3 vdd gnd cell_6t
Xbit_r4_c74 bl_74 br_74 wl_4 vdd gnd cell_6t
Xbit_r5_c74 bl_74 br_74 wl_5 vdd gnd cell_6t
Xbit_r6_c74 bl_74 br_74 wl_6 vdd gnd cell_6t
Xbit_r7_c74 bl_74 br_74 wl_7 vdd gnd cell_6t
Xbit_r8_c74 bl_74 br_74 wl_8 vdd gnd cell_6t
Xbit_r9_c74 bl_74 br_74 wl_9 vdd gnd cell_6t
Xbit_r10_c74 bl_74 br_74 wl_10 vdd gnd cell_6t
Xbit_r11_c74 bl_74 br_74 wl_11 vdd gnd cell_6t
Xbit_r12_c74 bl_74 br_74 wl_12 vdd gnd cell_6t
Xbit_r13_c74 bl_74 br_74 wl_13 vdd gnd cell_6t
Xbit_r14_c74 bl_74 br_74 wl_14 vdd gnd cell_6t
Xbit_r15_c74 bl_74 br_74 wl_15 vdd gnd cell_6t
Xbit_r16_c74 bl_74 br_74 wl_16 vdd gnd cell_6t
Xbit_r17_c74 bl_74 br_74 wl_17 vdd gnd cell_6t
Xbit_r18_c74 bl_74 br_74 wl_18 vdd gnd cell_6t
Xbit_r19_c74 bl_74 br_74 wl_19 vdd gnd cell_6t
Xbit_r20_c74 bl_74 br_74 wl_20 vdd gnd cell_6t
Xbit_r21_c74 bl_74 br_74 wl_21 vdd gnd cell_6t
Xbit_r22_c74 bl_74 br_74 wl_22 vdd gnd cell_6t
Xbit_r23_c74 bl_74 br_74 wl_23 vdd gnd cell_6t
Xbit_r24_c74 bl_74 br_74 wl_24 vdd gnd cell_6t
Xbit_r25_c74 bl_74 br_74 wl_25 vdd gnd cell_6t
Xbit_r26_c74 bl_74 br_74 wl_26 vdd gnd cell_6t
Xbit_r27_c74 bl_74 br_74 wl_27 vdd gnd cell_6t
Xbit_r28_c74 bl_74 br_74 wl_28 vdd gnd cell_6t
Xbit_r29_c74 bl_74 br_74 wl_29 vdd gnd cell_6t
Xbit_r30_c74 bl_74 br_74 wl_30 vdd gnd cell_6t
Xbit_r31_c74 bl_74 br_74 wl_31 vdd gnd cell_6t
Xbit_r32_c74 bl_74 br_74 wl_32 vdd gnd cell_6t
Xbit_r33_c74 bl_74 br_74 wl_33 vdd gnd cell_6t
Xbit_r34_c74 bl_74 br_74 wl_34 vdd gnd cell_6t
Xbit_r35_c74 bl_74 br_74 wl_35 vdd gnd cell_6t
Xbit_r36_c74 bl_74 br_74 wl_36 vdd gnd cell_6t
Xbit_r37_c74 bl_74 br_74 wl_37 vdd gnd cell_6t
Xbit_r38_c74 bl_74 br_74 wl_38 vdd gnd cell_6t
Xbit_r39_c74 bl_74 br_74 wl_39 vdd gnd cell_6t
Xbit_r40_c74 bl_74 br_74 wl_40 vdd gnd cell_6t
Xbit_r41_c74 bl_74 br_74 wl_41 vdd gnd cell_6t
Xbit_r42_c74 bl_74 br_74 wl_42 vdd gnd cell_6t
Xbit_r43_c74 bl_74 br_74 wl_43 vdd gnd cell_6t
Xbit_r44_c74 bl_74 br_74 wl_44 vdd gnd cell_6t
Xbit_r45_c74 bl_74 br_74 wl_45 vdd gnd cell_6t
Xbit_r46_c74 bl_74 br_74 wl_46 vdd gnd cell_6t
Xbit_r47_c74 bl_74 br_74 wl_47 vdd gnd cell_6t
Xbit_r48_c74 bl_74 br_74 wl_48 vdd gnd cell_6t
Xbit_r49_c74 bl_74 br_74 wl_49 vdd gnd cell_6t
Xbit_r50_c74 bl_74 br_74 wl_50 vdd gnd cell_6t
Xbit_r51_c74 bl_74 br_74 wl_51 vdd gnd cell_6t
Xbit_r52_c74 bl_74 br_74 wl_52 vdd gnd cell_6t
Xbit_r53_c74 bl_74 br_74 wl_53 vdd gnd cell_6t
Xbit_r54_c74 bl_74 br_74 wl_54 vdd gnd cell_6t
Xbit_r55_c74 bl_74 br_74 wl_55 vdd gnd cell_6t
Xbit_r56_c74 bl_74 br_74 wl_56 vdd gnd cell_6t
Xbit_r57_c74 bl_74 br_74 wl_57 vdd gnd cell_6t
Xbit_r58_c74 bl_74 br_74 wl_58 vdd gnd cell_6t
Xbit_r59_c74 bl_74 br_74 wl_59 vdd gnd cell_6t
Xbit_r60_c74 bl_74 br_74 wl_60 vdd gnd cell_6t
Xbit_r61_c74 bl_74 br_74 wl_61 vdd gnd cell_6t
Xbit_r62_c74 bl_74 br_74 wl_62 vdd gnd cell_6t
Xbit_r63_c74 bl_74 br_74 wl_63 vdd gnd cell_6t
Xbit_r64_c74 bl_74 br_74 wl_64 vdd gnd cell_6t
Xbit_r65_c74 bl_74 br_74 wl_65 vdd gnd cell_6t
Xbit_r66_c74 bl_74 br_74 wl_66 vdd gnd cell_6t
Xbit_r67_c74 bl_74 br_74 wl_67 vdd gnd cell_6t
Xbit_r68_c74 bl_74 br_74 wl_68 vdd gnd cell_6t
Xbit_r69_c74 bl_74 br_74 wl_69 vdd gnd cell_6t
Xbit_r70_c74 bl_74 br_74 wl_70 vdd gnd cell_6t
Xbit_r71_c74 bl_74 br_74 wl_71 vdd gnd cell_6t
Xbit_r72_c74 bl_74 br_74 wl_72 vdd gnd cell_6t
Xbit_r73_c74 bl_74 br_74 wl_73 vdd gnd cell_6t
Xbit_r74_c74 bl_74 br_74 wl_74 vdd gnd cell_6t
Xbit_r75_c74 bl_74 br_74 wl_75 vdd gnd cell_6t
Xbit_r76_c74 bl_74 br_74 wl_76 vdd gnd cell_6t
Xbit_r77_c74 bl_74 br_74 wl_77 vdd gnd cell_6t
Xbit_r78_c74 bl_74 br_74 wl_78 vdd gnd cell_6t
Xbit_r79_c74 bl_74 br_74 wl_79 vdd gnd cell_6t
Xbit_r80_c74 bl_74 br_74 wl_80 vdd gnd cell_6t
Xbit_r81_c74 bl_74 br_74 wl_81 vdd gnd cell_6t
Xbit_r82_c74 bl_74 br_74 wl_82 vdd gnd cell_6t
Xbit_r83_c74 bl_74 br_74 wl_83 vdd gnd cell_6t
Xbit_r84_c74 bl_74 br_74 wl_84 vdd gnd cell_6t
Xbit_r85_c74 bl_74 br_74 wl_85 vdd gnd cell_6t
Xbit_r86_c74 bl_74 br_74 wl_86 vdd gnd cell_6t
Xbit_r87_c74 bl_74 br_74 wl_87 vdd gnd cell_6t
Xbit_r88_c74 bl_74 br_74 wl_88 vdd gnd cell_6t
Xbit_r89_c74 bl_74 br_74 wl_89 vdd gnd cell_6t
Xbit_r90_c74 bl_74 br_74 wl_90 vdd gnd cell_6t
Xbit_r91_c74 bl_74 br_74 wl_91 vdd gnd cell_6t
Xbit_r92_c74 bl_74 br_74 wl_92 vdd gnd cell_6t
Xbit_r93_c74 bl_74 br_74 wl_93 vdd gnd cell_6t
Xbit_r94_c74 bl_74 br_74 wl_94 vdd gnd cell_6t
Xbit_r95_c74 bl_74 br_74 wl_95 vdd gnd cell_6t
Xbit_r96_c74 bl_74 br_74 wl_96 vdd gnd cell_6t
Xbit_r97_c74 bl_74 br_74 wl_97 vdd gnd cell_6t
Xbit_r98_c74 bl_74 br_74 wl_98 vdd gnd cell_6t
Xbit_r99_c74 bl_74 br_74 wl_99 vdd gnd cell_6t
Xbit_r100_c74 bl_74 br_74 wl_100 vdd gnd cell_6t
Xbit_r101_c74 bl_74 br_74 wl_101 vdd gnd cell_6t
Xbit_r102_c74 bl_74 br_74 wl_102 vdd gnd cell_6t
Xbit_r103_c74 bl_74 br_74 wl_103 vdd gnd cell_6t
Xbit_r104_c74 bl_74 br_74 wl_104 vdd gnd cell_6t
Xbit_r105_c74 bl_74 br_74 wl_105 vdd gnd cell_6t
Xbit_r106_c74 bl_74 br_74 wl_106 vdd gnd cell_6t
Xbit_r107_c74 bl_74 br_74 wl_107 vdd gnd cell_6t
Xbit_r108_c74 bl_74 br_74 wl_108 vdd gnd cell_6t
Xbit_r109_c74 bl_74 br_74 wl_109 vdd gnd cell_6t
Xbit_r110_c74 bl_74 br_74 wl_110 vdd gnd cell_6t
Xbit_r111_c74 bl_74 br_74 wl_111 vdd gnd cell_6t
Xbit_r112_c74 bl_74 br_74 wl_112 vdd gnd cell_6t
Xbit_r113_c74 bl_74 br_74 wl_113 vdd gnd cell_6t
Xbit_r114_c74 bl_74 br_74 wl_114 vdd gnd cell_6t
Xbit_r115_c74 bl_74 br_74 wl_115 vdd gnd cell_6t
Xbit_r116_c74 bl_74 br_74 wl_116 vdd gnd cell_6t
Xbit_r117_c74 bl_74 br_74 wl_117 vdd gnd cell_6t
Xbit_r118_c74 bl_74 br_74 wl_118 vdd gnd cell_6t
Xbit_r119_c74 bl_74 br_74 wl_119 vdd gnd cell_6t
Xbit_r120_c74 bl_74 br_74 wl_120 vdd gnd cell_6t
Xbit_r121_c74 bl_74 br_74 wl_121 vdd gnd cell_6t
Xbit_r122_c74 bl_74 br_74 wl_122 vdd gnd cell_6t
Xbit_r123_c74 bl_74 br_74 wl_123 vdd gnd cell_6t
Xbit_r124_c74 bl_74 br_74 wl_124 vdd gnd cell_6t
Xbit_r125_c74 bl_74 br_74 wl_125 vdd gnd cell_6t
Xbit_r126_c74 bl_74 br_74 wl_126 vdd gnd cell_6t
Xbit_r127_c74 bl_74 br_74 wl_127 vdd gnd cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd cell_6t
Xbit_r1_c75 bl_75 br_75 wl_1 vdd gnd cell_6t
Xbit_r2_c75 bl_75 br_75 wl_2 vdd gnd cell_6t
Xbit_r3_c75 bl_75 br_75 wl_3 vdd gnd cell_6t
Xbit_r4_c75 bl_75 br_75 wl_4 vdd gnd cell_6t
Xbit_r5_c75 bl_75 br_75 wl_5 vdd gnd cell_6t
Xbit_r6_c75 bl_75 br_75 wl_6 vdd gnd cell_6t
Xbit_r7_c75 bl_75 br_75 wl_7 vdd gnd cell_6t
Xbit_r8_c75 bl_75 br_75 wl_8 vdd gnd cell_6t
Xbit_r9_c75 bl_75 br_75 wl_9 vdd gnd cell_6t
Xbit_r10_c75 bl_75 br_75 wl_10 vdd gnd cell_6t
Xbit_r11_c75 bl_75 br_75 wl_11 vdd gnd cell_6t
Xbit_r12_c75 bl_75 br_75 wl_12 vdd gnd cell_6t
Xbit_r13_c75 bl_75 br_75 wl_13 vdd gnd cell_6t
Xbit_r14_c75 bl_75 br_75 wl_14 vdd gnd cell_6t
Xbit_r15_c75 bl_75 br_75 wl_15 vdd gnd cell_6t
Xbit_r16_c75 bl_75 br_75 wl_16 vdd gnd cell_6t
Xbit_r17_c75 bl_75 br_75 wl_17 vdd gnd cell_6t
Xbit_r18_c75 bl_75 br_75 wl_18 vdd gnd cell_6t
Xbit_r19_c75 bl_75 br_75 wl_19 vdd gnd cell_6t
Xbit_r20_c75 bl_75 br_75 wl_20 vdd gnd cell_6t
Xbit_r21_c75 bl_75 br_75 wl_21 vdd gnd cell_6t
Xbit_r22_c75 bl_75 br_75 wl_22 vdd gnd cell_6t
Xbit_r23_c75 bl_75 br_75 wl_23 vdd gnd cell_6t
Xbit_r24_c75 bl_75 br_75 wl_24 vdd gnd cell_6t
Xbit_r25_c75 bl_75 br_75 wl_25 vdd gnd cell_6t
Xbit_r26_c75 bl_75 br_75 wl_26 vdd gnd cell_6t
Xbit_r27_c75 bl_75 br_75 wl_27 vdd gnd cell_6t
Xbit_r28_c75 bl_75 br_75 wl_28 vdd gnd cell_6t
Xbit_r29_c75 bl_75 br_75 wl_29 vdd gnd cell_6t
Xbit_r30_c75 bl_75 br_75 wl_30 vdd gnd cell_6t
Xbit_r31_c75 bl_75 br_75 wl_31 vdd gnd cell_6t
Xbit_r32_c75 bl_75 br_75 wl_32 vdd gnd cell_6t
Xbit_r33_c75 bl_75 br_75 wl_33 vdd gnd cell_6t
Xbit_r34_c75 bl_75 br_75 wl_34 vdd gnd cell_6t
Xbit_r35_c75 bl_75 br_75 wl_35 vdd gnd cell_6t
Xbit_r36_c75 bl_75 br_75 wl_36 vdd gnd cell_6t
Xbit_r37_c75 bl_75 br_75 wl_37 vdd gnd cell_6t
Xbit_r38_c75 bl_75 br_75 wl_38 vdd gnd cell_6t
Xbit_r39_c75 bl_75 br_75 wl_39 vdd gnd cell_6t
Xbit_r40_c75 bl_75 br_75 wl_40 vdd gnd cell_6t
Xbit_r41_c75 bl_75 br_75 wl_41 vdd gnd cell_6t
Xbit_r42_c75 bl_75 br_75 wl_42 vdd gnd cell_6t
Xbit_r43_c75 bl_75 br_75 wl_43 vdd gnd cell_6t
Xbit_r44_c75 bl_75 br_75 wl_44 vdd gnd cell_6t
Xbit_r45_c75 bl_75 br_75 wl_45 vdd gnd cell_6t
Xbit_r46_c75 bl_75 br_75 wl_46 vdd gnd cell_6t
Xbit_r47_c75 bl_75 br_75 wl_47 vdd gnd cell_6t
Xbit_r48_c75 bl_75 br_75 wl_48 vdd gnd cell_6t
Xbit_r49_c75 bl_75 br_75 wl_49 vdd gnd cell_6t
Xbit_r50_c75 bl_75 br_75 wl_50 vdd gnd cell_6t
Xbit_r51_c75 bl_75 br_75 wl_51 vdd gnd cell_6t
Xbit_r52_c75 bl_75 br_75 wl_52 vdd gnd cell_6t
Xbit_r53_c75 bl_75 br_75 wl_53 vdd gnd cell_6t
Xbit_r54_c75 bl_75 br_75 wl_54 vdd gnd cell_6t
Xbit_r55_c75 bl_75 br_75 wl_55 vdd gnd cell_6t
Xbit_r56_c75 bl_75 br_75 wl_56 vdd gnd cell_6t
Xbit_r57_c75 bl_75 br_75 wl_57 vdd gnd cell_6t
Xbit_r58_c75 bl_75 br_75 wl_58 vdd gnd cell_6t
Xbit_r59_c75 bl_75 br_75 wl_59 vdd gnd cell_6t
Xbit_r60_c75 bl_75 br_75 wl_60 vdd gnd cell_6t
Xbit_r61_c75 bl_75 br_75 wl_61 vdd gnd cell_6t
Xbit_r62_c75 bl_75 br_75 wl_62 vdd gnd cell_6t
Xbit_r63_c75 bl_75 br_75 wl_63 vdd gnd cell_6t
Xbit_r64_c75 bl_75 br_75 wl_64 vdd gnd cell_6t
Xbit_r65_c75 bl_75 br_75 wl_65 vdd gnd cell_6t
Xbit_r66_c75 bl_75 br_75 wl_66 vdd gnd cell_6t
Xbit_r67_c75 bl_75 br_75 wl_67 vdd gnd cell_6t
Xbit_r68_c75 bl_75 br_75 wl_68 vdd gnd cell_6t
Xbit_r69_c75 bl_75 br_75 wl_69 vdd gnd cell_6t
Xbit_r70_c75 bl_75 br_75 wl_70 vdd gnd cell_6t
Xbit_r71_c75 bl_75 br_75 wl_71 vdd gnd cell_6t
Xbit_r72_c75 bl_75 br_75 wl_72 vdd gnd cell_6t
Xbit_r73_c75 bl_75 br_75 wl_73 vdd gnd cell_6t
Xbit_r74_c75 bl_75 br_75 wl_74 vdd gnd cell_6t
Xbit_r75_c75 bl_75 br_75 wl_75 vdd gnd cell_6t
Xbit_r76_c75 bl_75 br_75 wl_76 vdd gnd cell_6t
Xbit_r77_c75 bl_75 br_75 wl_77 vdd gnd cell_6t
Xbit_r78_c75 bl_75 br_75 wl_78 vdd gnd cell_6t
Xbit_r79_c75 bl_75 br_75 wl_79 vdd gnd cell_6t
Xbit_r80_c75 bl_75 br_75 wl_80 vdd gnd cell_6t
Xbit_r81_c75 bl_75 br_75 wl_81 vdd gnd cell_6t
Xbit_r82_c75 bl_75 br_75 wl_82 vdd gnd cell_6t
Xbit_r83_c75 bl_75 br_75 wl_83 vdd gnd cell_6t
Xbit_r84_c75 bl_75 br_75 wl_84 vdd gnd cell_6t
Xbit_r85_c75 bl_75 br_75 wl_85 vdd gnd cell_6t
Xbit_r86_c75 bl_75 br_75 wl_86 vdd gnd cell_6t
Xbit_r87_c75 bl_75 br_75 wl_87 vdd gnd cell_6t
Xbit_r88_c75 bl_75 br_75 wl_88 vdd gnd cell_6t
Xbit_r89_c75 bl_75 br_75 wl_89 vdd gnd cell_6t
Xbit_r90_c75 bl_75 br_75 wl_90 vdd gnd cell_6t
Xbit_r91_c75 bl_75 br_75 wl_91 vdd gnd cell_6t
Xbit_r92_c75 bl_75 br_75 wl_92 vdd gnd cell_6t
Xbit_r93_c75 bl_75 br_75 wl_93 vdd gnd cell_6t
Xbit_r94_c75 bl_75 br_75 wl_94 vdd gnd cell_6t
Xbit_r95_c75 bl_75 br_75 wl_95 vdd gnd cell_6t
Xbit_r96_c75 bl_75 br_75 wl_96 vdd gnd cell_6t
Xbit_r97_c75 bl_75 br_75 wl_97 vdd gnd cell_6t
Xbit_r98_c75 bl_75 br_75 wl_98 vdd gnd cell_6t
Xbit_r99_c75 bl_75 br_75 wl_99 vdd gnd cell_6t
Xbit_r100_c75 bl_75 br_75 wl_100 vdd gnd cell_6t
Xbit_r101_c75 bl_75 br_75 wl_101 vdd gnd cell_6t
Xbit_r102_c75 bl_75 br_75 wl_102 vdd gnd cell_6t
Xbit_r103_c75 bl_75 br_75 wl_103 vdd gnd cell_6t
Xbit_r104_c75 bl_75 br_75 wl_104 vdd gnd cell_6t
Xbit_r105_c75 bl_75 br_75 wl_105 vdd gnd cell_6t
Xbit_r106_c75 bl_75 br_75 wl_106 vdd gnd cell_6t
Xbit_r107_c75 bl_75 br_75 wl_107 vdd gnd cell_6t
Xbit_r108_c75 bl_75 br_75 wl_108 vdd gnd cell_6t
Xbit_r109_c75 bl_75 br_75 wl_109 vdd gnd cell_6t
Xbit_r110_c75 bl_75 br_75 wl_110 vdd gnd cell_6t
Xbit_r111_c75 bl_75 br_75 wl_111 vdd gnd cell_6t
Xbit_r112_c75 bl_75 br_75 wl_112 vdd gnd cell_6t
Xbit_r113_c75 bl_75 br_75 wl_113 vdd gnd cell_6t
Xbit_r114_c75 bl_75 br_75 wl_114 vdd gnd cell_6t
Xbit_r115_c75 bl_75 br_75 wl_115 vdd gnd cell_6t
Xbit_r116_c75 bl_75 br_75 wl_116 vdd gnd cell_6t
Xbit_r117_c75 bl_75 br_75 wl_117 vdd gnd cell_6t
Xbit_r118_c75 bl_75 br_75 wl_118 vdd gnd cell_6t
Xbit_r119_c75 bl_75 br_75 wl_119 vdd gnd cell_6t
Xbit_r120_c75 bl_75 br_75 wl_120 vdd gnd cell_6t
Xbit_r121_c75 bl_75 br_75 wl_121 vdd gnd cell_6t
Xbit_r122_c75 bl_75 br_75 wl_122 vdd gnd cell_6t
Xbit_r123_c75 bl_75 br_75 wl_123 vdd gnd cell_6t
Xbit_r124_c75 bl_75 br_75 wl_124 vdd gnd cell_6t
Xbit_r125_c75 bl_75 br_75 wl_125 vdd gnd cell_6t
Xbit_r126_c75 bl_75 br_75 wl_126 vdd gnd cell_6t
Xbit_r127_c75 bl_75 br_75 wl_127 vdd gnd cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd cell_6t
Xbit_r1_c76 bl_76 br_76 wl_1 vdd gnd cell_6t
Xbit_r2_c76 bl_76 br_76 wl_2 vdd gnd cell_6t
Xbit_r3_c76 bl_76 br_76 wl_3 vdd gnd cell_6t
Xbit_r4_c76 bl_76 br_76 wl_4 vdd gnd cell_6t
Xbit_r5_c76 bl_76 br_76 wl_5 vdd gnd cell_6t
Xbit_r6_c76 bl_76 br_76 wl_6 vdd gnd cell_6t
Xbit_r7_c76 bl_76 br_76 wl_7 vdd gnd cell_6t
Xbit_r8_c76 bl_76 br_76 wl_8 vdd gnd cell_6t
Xbit_r9_c76 bl_76 br_76 wl_9 vdd gnd cell_6t
Xbit_r10_c76 bl_76 br_76 wl_10 vdd gnd cell_6t
Xbit_r11_c76 bl_76 br_76 wl_11 vdd gnd cell_6t
Xbit_r12_c76 bl_76 br_76 wl_12 vdd gnd cell_6t
Xbit_r13_c76 bl_76 br_76 wl_13 vdd gnd cell_6t
Xbit_r14_c76 bl_76 br_76 wl_14 vdd gnd cell_6t
Xbit_r15_c76 bl_76 br_76 wl_15 vdd gnd cell_6t
Xbit_r16_c76 bl_76 br_76 wl_16 vdd gnd cell_6t
Xbit_r17_c76 bl_76 br_76 wl_17 vdd gnd cell_6t
Xbit_r18_c76 bl_76 br_76 wl_18 vdd gnd cell_6t
Xbit_r19_c76 bl_76 br_76 wl_19 vdd gnd cell_6t
Xbit_r20_c76 bl_76 br_76 wl_20 vdd gnd cell_6t
Xbit_r21_c76 bl_76 br_76 wl_21 vdd gnd cell_6t
Xbit_r22_c76 bl_76 br_76 wl_22 vdd gnd cell_6t
Xbit_r23_c76 bl_76 br_76 wl_23 vdd gnd cell_6t
Xbit_r24_c76 bl_76 br_76 wl_24 vdd gnd cell_6t
Xbit_r25_c76 bl_76 br_76 wl_25 vdd gnd cell_6t
Xbit_r26_c76 bl_76 br_76 wl_26 vdd gnd cell_6t
Xbit_r27_c76 bl_76 br_76 wl_27 vdd gnd cell_6t
Xbit_r28_c76 bl_76 br_76 wl_28 vdd gnd cell_6t
Xbit_r29_c76 bl_76 br_76 wl_29 vdd gnd cell_6t
Xbit_r30_c76 bl_76 br_76 wl_30 vdd gnd cell_6t
Xbit_r31_c76 bl_76 br_76 wl_31 vdd gnd cell_6t
Xbit_r32_c76 bl_76 br_76 wl_32 vdd gnd cell_6t
Xbit_r33_c76 bl_76 br_76 wl_33 vdd gnd cell_6t
Xbit_r34_c76 bl_76 br_76 wl_34 vdd gnd cell_6t
Xbit_r35_c76 bl_76 br_76 wl_35 vdd gnd cell_6t
Xbit_r36_c76 bl_76 br_76 wl_36 vdd gnd cell_6t
Xbit_r37_c76 bl_76 br_76 wl_37 vdd gnd cell_6t
Xbit_r38_c76 bl_76 br_76 wl_38 vdd gnd cell_6t
Xbit_r39_c76 bl_76 br_76 wl_39 vdd gnd cell_6t
Xbit_r40_c76 bl_76 br_76 wl_40 vdd gnd cell_6t
Xbit_r41_c76 bl_76 br_76 wl_41 vdd gnd cell_6t
Xbit_r42_c76 bl_76 br_76 wl_42 vdd gnd cell_6t
Xbit_r43_c76 bl_76 br_76 wl_43 vdd gnd cell_6t
Xbit_r44_c76 bl_76 br_76 wl_44 vdd gnd cell_6t
Xbit_r45_c76 bl_76 br_76 wl_45 vdd gnd cell_6t
Xbit_r46_c76 bl_76 br_76 wl_46 vdd gnd cell_6t
Xbit_r47_c76 bl_76 br_76 wl_47 vdd gnd cell_6t
Xbit_r48_c76 bl_76 br_76 wl_48 vdd gnd cell_6t
Xbit_r49_c76 bl_76 br_76 wl_49 vdd gnd cell_6t
Xbit_r50_c76 bl_76 br_76 wl_50 vdd gnd cell_6t
Xbit_r51_c76 bl_76 br_76 wl_51 vdd gnd cell_6t
Xbit_r52_c76 bl_76 br_76 wl_52 vdd gnd cell_6t
Xbit_r53_c76 bl_76 br_76 wl_53 vdd gnd cell_6t
Xbit_r54_c76 bl_76 br_76 wl_54 vdd gnd cell_6t
Xbit_r55_c76 bl_76 br_76 wl_55 vdd gnd cell_6t
Xbit_r56_c76 bl_76 br_76 wl_56 vdd gnd cell_6t
Xbit_r57_c76 bl_76 br_76 wl_57 vdd gnd cell_6t
Xbit_r58_c76 bl_76 br_76 wl_58 vdd gnd cell_6t
Xbit_r59_c76 bl_76 br_76 wl_59 vdd gnd cell_6t
Xbit_r60_c76 bl_76 br_76 wl_60 vdd gnd cell_6t
Xbit_r61_c76 bl_76 br_76 wl_61 vdd gnd cell_6t
Xbit_r62_c76 bl_76 br_76 wl_62 vdd gnd cell_6t
Xbit_r63_c76 bl_76 br_76 wl_63 vdd gnd cell_6t
Xbit_r64_c76 bl_76 br_76 wl_64 vdd gnd cell_6t
Xbit_r65_c76 bl_76 br_76 wl_65 vdd gnd cell_6t
Xbit_r66_c76 bl_76 br_76 wl_66 vdd gnd cell_6t
Xbit_r67_c76 bl_76 br_76 wl_67 vdd gnd cell_6t
Xbit_r68_c76 bl_76 br_76 wl_68 vdd gnd cell_6t
Xbit_r69_c76 bl_76 br_76 wl_69 vdd gnd cell_6t
Xbit_r70_c76 bl_76 br_76 wl_70 vdd gnd cell_6t
Xbit_r71_c76 bl_76 br_76 wl_71 vdd gnd cell_6t
Xbit_r72_c76 bl_76 br_76 wl_72 vdd gnd cell_6t
Xbit_r73_c76 bl_76 br_76 wl_73 vdd gnd cell_6t
Xbit_r74_c76 bl_76 br_76 wl_74 vdd gnd cell_6t
Xbit_r75_c76 bl_76 br_76 wl_75 vdd gnd cell_6t
Xbit_r76_c76 bl_76 br_76 wl_76 vdd gnd cell_6t
Xbit_r77_c76 bl_76 br_76 wl_77 vdd gnd cell_6t
Xbit_r78_c76 bl_76 br_76 wl_78 vdd gnd cell_6t
Xbit_r79_c76 bl_76 br_76 wl_79 vdd gnd cell_6t
Xbit_r80_c76 bl_76 br_76 wl_80 vdd gnd cell_6t
Xbit_r81_c76 bl_76 br_76 wl_81 vdd gnd cell_6t
Xbit_r82_c76 bl_76 br_76 wl_82 vdd gnd cell_6t
Xbit_r83_c76 bl_76 br_76 wl_83 vdd gnd cell_6t
Xbit_r84_c76 bl_76 br_76 wl_84 vdd gnd cell_6t
Xbit_r85_c76 bl_76 br_76 wl_85 vdd gnd cell_6t
Xbit_r86_c76 bl_76 br_76 wl_86 vdd gnd cell_6t
Xbit_r87_c76 bl_76 br_76 wl_87 vdd gnd cell_6t
Xbit_r88_c76 bl_76 br_76 wl_88 vdd gnd cell_6t
Xbit_r89_c76 bl_76 br_76 wl_89 vdd gnd cell_6t
Xbit_r90_c76 bl_76 br_76 wl_90 vdd gnd cell_6t
Xbit_r91_c76 bl_76 br_76 wl_91 vdd gnd cell_6t
Xbit_r92_c76 bl_76 br_76 wl_92 vdd gnd cell_6t
Xbit_r93_c76 bl_76 br_76 wl_93 vdd gnd cell_6t
Xbit_r94_c76 bl_76 br_76 wl_94 vdd gnd cell_6t
Xbit_r95_c76 bl_76 br_76 wl_95 vdd gnd cell_6t
Xbit_r96_c76 bl_76 br_76 wl_96 vdd gnd cell_6t
Xbit_r97_c76 bl_76 br_76 wl_97 vdd gnd cell_6t
Xbit_r98_c76 bl_76 br_76 wl_98 vdd gnd cell_6t
Xbit_r99_c76 bl_76 br_76 wl_99 vdd gnd cell_6t
Xbit_r100_c76 bl_76 br_76 wl_100 vdd gnd cell_6t
Xbit_r101_c76 bl_76 br_76 wl_101 vdd gnd cell_6t
Xbit_r102_c76 bl_76 br_76 wl_102 vdd gnd cell_6t
Xbit_r103_c76 bl_76 br_76 wl_103 vdd gnd cell_6t
Xbit_r104_c76 bl_76 br_76 wl_104 vdd gnd cell_6t
Xbit_r105_c76 bl_76 br_76 wl_105 vdd gnd cell_6t
Xbit_r106_c76 bl_76 br_76 wl_106 vdd gnd cell_6t
Xbit_r107_c76 bl_76 br_76 wl_107 vdd gnd cell_6t
Xbit_r108_c76 bl_76 br_76 wl_108 vdd gnd cell_6t
Xbit_r109_c76 bl_76 br_76 wl_109 vdd gnd cell_6t
Xbit_r110_c76 bl_76 br_76 wl_110 vdd gnd cell_6t
Xbit_r111_c76 bl_76 br_76 wl_111 vdd gnd cell_6t
Xbit_r112_c76 bl_76 br_76 wl_112 vdd gnd cell_6t
Xbit_r113_c76 bl_76 br_76 wl_113 vdd gnd cell_6t
Xbit_r114_c76 bl_76 br_76 wl_114 vdd gnd cell_6t
Xbit_r115_c76 bl_76 br_76 wl_115 vdd gnd cell_6t
Xbit_r116_c76 bl_76 br_76 wl_116 vdd gnd cell_6t
Xbit_r117_c76 bl_76 br_76 wl_117 vdd gnd cell_6t
Xbit_r118_c76 bl_76 br_76 wl_118 vdd gnd cell_6t
Xbit_r119_c76 bl_76 br_76 wl_119 vdd gnd cell_6t
Xbit_r120_c76 bl_76 br_76 wl_120 vdd gnd cell_6t
Xbit_r121_c76 bl_76 br_76 wl_121 vdd gnd cell_6t
Xbit_r122_c76 bl_76 br_76 wl_122 vdd gnd cell_6t
Xbit_r123_c76 bl_76 br_76 wl_123 vdd gnd cell_6t
Xbit_r124_c76 bl_76 br_76 wl_124 vdd gnd cell_6t
Xbit_r125_c76 bl_76 br_76 wl_125 vdd gnd cell_6t
Xbit_r126_c76 bl_76 br_76 wl_126 vdd gnd cell_6t
Xbit_r127_c76 bl_76 br_76 wl_127 vdd gnd cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd cell_6t
Xbit_r1_c77 bl_77 br_77 wl_1 vdd gnd cell_6t
Xbit_r2_c77 bl_77 br_77 wl_2 vdd gnd cell_6t
Xbit_r3_c77 bl_77 br_77 wl_3 vdd gnd cell_6t
Xbit_r4_c77 bl_77 br_77 wl_4 vdd gnd cell_6t
Xbit_r5_c77 bl_77 br_77 wl_5 vdd gnd cell_6t
Xbit_r6_c77 bl_77 br_77 wl_6 vdd gnd cell_6t
Xbit_r7_c77 bl_77 br_77 wl_7 vdd gnd cell_6t
Xbit_r8_c77 bl_77 br_77 wl_8 vdd gnd cell_6t
Xbit_r9_c77 bl_77 br_77 wl_9 vdd gnd cell_6t
Xbit_r10_c77 bl_77 br_77 wl_10 vdd gnd cell_6t
Xbit_r11_c77 bl_77 br_77 wl_11 vdd gnd cell_6t
Xbit_r12_c77 bl_77 br_77 wl_12 vdd gnd cell_6t
Xbit_r13_c77 bl_77 br_77 wl_13 vdd gnd cell_6t
Xbit_r14_c77 bl_77 br_77 wl_14 vdd gnd cell_6t
Xbit_r15_c77 bl_77 br_77 wl_15 vdd gnd cell_6t
Xbit_r16_c77 bl_77 br_77 wl_16 vdd gnd cell_6t
Xbit_r17_c77 bl_77 br_77 wl_17 vdd gnd cell_6t
Xbit_r18_c77 bl_77 br_77 wl_18 vdd gnd cell_6t
Xbit_r19_c77 bl_77 br_77 wl_19 vdd gnd cell_6t
Xbit_r20_c77 bl_77 br_77 wl_20 vdd gnd cell_6t
Xbit_r21_c77 bl_77 br_77 wl_21 vdd gnd cell_6t
Xbit_r22_c77 bl_77 br_77 wl_22 vdd gnd cell_6t
Xbit_r23_c77 bl_77 br_77 wl_23 vdd gnd cell_6t
Xbit_r24_c77 bl_77 br_77 wl_24 vdd gnd cell_6t
Xbit_r25_c77 bl_77 br_77 wl_25 vdd gnd cell_6t
Xbit_r26_c77 bl_77 br_77 wl_26 vdd gnd cell_6t
Xbit_r27_c77 bl_77 br_77 wl_27 vdd gnd cell_6t
Xbit_r28_c77 bl_77 br_77 wl_28 vdd gnd cell_6t
Xbit_r29_c77 bl_77 br_77 wl_29 vdd gnd cell_6t
Xbit_r30_c77 bl_77 br_77 wl_30 vdd gnd cell_6t
Xbit_r31_c77 bl_77 br_77 wl_31 vdd gnd cell_6t
Xbit_r32_c77 bl_77 br_77 wl_32 vdd gnd cell_6t
Xbit_r33_c77 bl_77 br_77 wl_33 vdd gnd cell_6t
Xbit_r34_c77 bl_77 br_77 wl_34 vdd gnd cell_6t
Xbit_r35_c77 bl_77 br_77 wl_35 vdd gnd cell_6t
Xbit_r36_c77 bl_77 br_77 wl_36 vdd gnd cell_6t
Xbit_r37_c77 bl_77 br_77 wl_37 vdd gnd cell_6t
Xbit_r38_c77 bl_77 br_77 wl_38 vdd gnd cell_6t
Xbit_r39_c77 bl_77 br_77 wl_39 vdd gnd cell_6t
Xbit_r40_c77 bl_77 br_77 wl_40 vdd gnd cell_6t
Xbit_r41_c77 bl_77 br_77 wl_41 vdd gnd cell_6t
Xbit_r42_c77 bl_77 br_77 wl_42 vdd gnd cell_6t
Xbit_r43_c77 bl_77 br_77 wl_43 vdd gnd cell_6t
Xbit_r44_c77 bl_77 br_77 wl_44 vdd gnd cell_6t
Xbit_r45_c77 bl_77 br_77 wl_45 vdd gnd cell_6t
Xbit_r46_c77 bl_77 br_77 wl_46 vdd gnd cell_6t
Xbit_r47_c77 bl_77 br_77 wl_47 vdd gnd cell_6t
Xbit_r48_c77 bl_77 br_77 wl_48 vdd gnd cell_6t
Xbit_r49_c77 bl_77 br_77 wl_49 vdd gnd cell_6t
Xbit_r50_c77 bl_77 br_77 wl_50 vdd gnd cell_6t
Xbit_r51_c77 bl_77 br_77 wl_51 vdd gnd cell_6t
Xbit_r52_c77 bl_77 br_77 wl_52 vdd gnd cell_6t
Xbit_r53_c77 bl_77 br_77 wl_53 vdd gnd cell_6t
Xbit_r54_c77 bl_77 br_77 wl_54 vdd gnd cell_6t
Xbit_r55_c77 bl_77 br_77 wl_55 vdd gnd cell_6t
Xbit_r56_c77 bl_77 br_77 wl_56 vdd gnd cell_6t
Xbit_r57_c77 bl_77 br_77 wl_57 vdd gnd cell_6t
Xbit_r58_c77 bl_77 br_77 wl_58 vdd gnd cell_6t
Xbit_r59_c77 bl_77 br_77 wl_59 vdd gnd cell_6t
Xbit_r60_c77 bl_77 br_77 wl_60 vdd gnd cell_6t
Xbit_r61_c77 bl_77 br_77 wl_61 vdd gnd cell_6t
Xbit_r62_c77 bl_77 br_77 wl_62 vdd gnd cell_6t
Xbit_r63_c77 bl_77 br_77 wl_63 vdd gnd cell_6t
Xbit_r64_c77 bl_77 br_77 wl_64 vdd gnd cell_6t
Xbit_r65_c77 bl_77 br_77 wl_65 vdd gnd cell_6t
Xbit_r66_c77 bl_77 br_77 wl_66 vdd gnd cell_6t
Xbit_r67_c77 bl_77 br_77 wl_67 vdd gnd cell_6t
Xbit_r68_c77 bl_77 br_77 wl_68 vdd gnd cell_6t
Xbit_r69_c77 bl_77 br_77 wl_69 vdd gnd cell_6t
Xbit_r70_c77 bl_77 br_77 wl_70 vdd gnd cell_6t
Xbit_r71_c77 bl_77 br_77 wl_71 vdd gnd cell_6t
Xbit_r72_c77 bl_77 br_77 wl_72 vdd gnd cell_6t
Xbit_r73_c77 bl_77 br_77 wl_73 vdd gnd cell_6t
Xbit_r74_c77 bl_77 br_77 wl_74 vdd gnd cell_6t
Xbit_r75_c77 bl_77 br_77 wl_75 vdd gnd cell_6t
Xbit_r76_c77 bl_77 br_77 wl_76 vdd gnd cell_6t
Xbit_r77_c77 bl_77 br_77 wl_77 vdd gnd cell_6t
Xbit_r78_c77 bl_77 br_77 wl_78 vdd gnd cell_6t
Xbit_r79_c77 bl_77 br_77 wl_79 vdd gnd cell_6t
Xbit_r80_c77 bl_77 br_77 wl_80 vdd gnd cell_6t
Xbit_r81_c77 bl_77 br_77 wl_81 vdd gnd cell_6t
Xbit_r82_c77 bl_77 br_77 wl_82 vdd gnd cell_6t
Xbit_r83_c77 bl_77 br_77 wl_83 vdd gnd cell_6t
Xbit_r84_c77 bl_77 br_77 wl_84 vdd gnd cell_6t
Xbit_r85_c77 bl_77 br_77 wl_85 vdd gnd cell_6t
Xbit_r86_c77 bl_77 br_77 wl_86 vdd gnd cell_6t
Xbit_r87_c77 bl_77 br_77 wl_87 vdd gnd cell_6t
Xbit_r88_c77 bl_77 br_77 wl_88 vdd gnd cell_6t
Xbit_r89_c77 bl_77 br_77 wl_89 vdd gnd cell_6t
Xbit_r90_c77 bl_77 br_77 wl_90 vdd gnd cell_6t
Xbit_r91_c77 bl_77 br_77 wl_91 vdd gnd cell_6t
Xbit_r92_c77 bl_77 br_77 wl_92 vdd gnd cell_6t
Xbit_r93_c77 bl_77 br_77 wl_93 vdd gnd cell_6t
Xbit_r94_c77 bl_77 br_77 wl_94 vdd gnd cell_6t
Xbit_r95_c77 bl_77 br_77 wl_95 vdd gnd cell_6t
Xbit_r96_c77 bl_77 br_77 wl_96 vdd gnd cell_6t
Xbit_r97_c77 bl_77 br_77 wl_97 vdd gnd cell_6t
Xbit_r98_c77 bl_77 br_77 wl_98 vdd gnd cell_6t
Xbit_r99_c77 bl_77 br_77 wl_99 vdd gnd cell_6t
Xbit_r100_c77 bl_77 br_77 wl_100 vdd gnd cell_6t
Xbit_r101_c77 bl_77 br_77 wl_101 vdd gnd cell_6t
Xbit_r102_c77 bl_77 br_77 wl_102 vdd gnd cell_6t
Xbit_r103_c77 bl_77 br_77 wl_103 vdd gnd cell_6t
Xbit_r104_c77 bl_77 br_77 wl_104 vdd gnd cell_6t
Xbit_r105_c77 bl_77 br_77 wl_105 vdd gnd cell_6t
Xbit_r106_c77 bl_77 br_77 wl_106 vdd gnd cell_6t
Xbit_r107_c77 bl_77 br_77 wl_107 vdd gnd cell_6t
Xbit_r108_c77 bl_77 br_77 wl_108 vdd gnd cell_6t
Xbit_r109_c77 bl_77 br_77 wl_109 vdd gnd cell_6t
Xbit_r110_c77 bl_77 br_77 wl_110 vdd gnd cell_6t
Xbit_r111_c77 bl_77 br_77 wl_111 vdd gnd cell_6t
Xbit_r112_c77 bl_77 br_77 wl_112 vdd gnd cell_6t
Xbit_r113_c77 bl_77 br_77 wl_113 vdd gnd cell_6t
Xbit_r114_c77 bl_77 br_77 wl_114 vdd gnd cell_6t
Xbit_r115_c77 bl_77 br_77 wl_115 vdd gnd cell_6t
Xbit_r116_c77 bl_77 br_77 wl_116 vdd gnd cell_6t
Xbit_r117_c77 bl_77 br_77 wl_117 vdd gnd cell_6t
Xbit_r118_c77 bl_77 br_77 wl_118 vdd gnd cell_6t
Xbit_r119_c77 bl_77 br_77 wl_119 vdd gnd cell_6t
Xbit_r120_c77 bl_77 br_77 wl_120 vdd gnd cell_6t
Xbit_r121_c77 bl_77 br_77 wl_121 vdd gnd cell_6t
Xbit_r122_c77 bl_77 br_77 wl_122 vdd gnd cell_6t
Xbit_r123_c77 bl_77 br_77 wl_123 vdd gnd cell_6t
Xbit_r124_c77 bl_77 br_77 wl_124 vdd gnd cell_6t
Xbit_r125_c77 bl_77 br_77 wl_125 vdd gnd cell_6t
Xbit_r126_c77 bl_77 br_77 wl_126 vdd gnd cell_6t
Xbit_r127_c77 bl_77 br_77 wl_127 vdd gnd cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd cell_6t
Xbit_r1_c78 bl_78 br_78 wl_1 vdd gnd cell_6t
Xbit_r2_c78 bl_78 br_78 wl_2 vdd gnd cell_6t
Xbit_r3_c78 bl_78 br_78 wl_3 vdd gnd cell_6t
Xbit_r4_c78 bl_78 br_78 wl_4 vdd gnd cell_6t
Xbit_r5_c78 bl_78 br_78 wl_5 vdd gnd cell_6t
Xbit_r6_c78 bl_78 br_78 wl_6 vdd gnd cell_6t
Xbit_r7_c78 bl_78 br_78 wl_7 vdd gnd cell_6t
Xbit_r8_c78 bl_78 br_78 wl_8 vdd gnd cell_6t
Xbit_r9_c78 bl_78 br_78 wl_9 vdd gnd cell_6t
Xbit_r10_c78 bl_78 br_78 wl_10 vdd gnd cell_6t
Xbit_r11_c78 bl_78 br_78 wl_11 vdd gnd cell_6t
Xbit_r12_c78 bl_78 br_78 wl_12 vdd gnd cell_6t
Xbit_r13_c78 bl_78 br_78 wl_13 vdd gnd cell_6t
Xbit_r14_c78 bl_78 br_78 wl_14 vdd gnd cell_6t
Xbit_r15_c78 bl_78 br_78 wl_15 vdd gnd cell_6t
Xbit_r16_c78 bl_78 br_78 wl_16 vdd gnd cell_6t
Xbit_r17_c78 bl_78 br_78 wl_17 vdd gnd cell_6t
Xbit_r18_c78 bl_78 br_78 wl_18 vdd gnd cell_6t
Xbit_r19_c78 bl_78 br_78 wl_19 vdd gnd cell_6t
Xbit_r20_c78 bl_78 br_78 wl_20 vdd gnd cell_6t
Xbit_r21_c78 bl_78 br_78 wl_21 vdd gnd cell_6t
Xbit_r22_c78 bl_78 br_78 wl_22 vdd gnd cell_6t
Xbit_r23_c78 bl_78 br_78 wl_23 vdd gnd cell_6t
Xbit_r24_c78 bl_78 br_78 wl_24 vdd gnd cell_6t
Xbit_r25_c78 bl_78 br_78 wl_25 vdd gnd cell_6t
Xbit_r26_c78 bl_78 br_78 wl_26 vdd gnd cell_6t
Xbit_r27_c78 bl_78 br_78 wl_27 vdd gnd cell_6t
Xbit_r28_c78 bl_78 br_78 wl_28 vdd gnd cell_6t
Xbit_r29_c78 bl_78 br_78 wl_29 vdd gnd cell_6t
Xbit_r30_c78 bl_78 br_78 wl_30 vdd gnd cell_6t
Xbit_r31_c78 bl_78 br_78 wl_31 vdd gnd cell_6t
Xbit_r32_c78 bl_78 br_78 wl_32 vdd gnd cell_6t
Xbit_r33_c78 bl_78 br_78 wl_33 vdd gnd cell_6t
Xbit_r34_c78 bl_78 br_78 wl_34 vdd gnd cell_6t
Xbit_r35_c78 bl_78 br_78 wl_35 vdd gnd cell_6t
Xbit_r36_c78 bl_78 br_78 wl_36 vdd gnd cell_6t
Xbit_r37_c78 bl_78 br_78 wl_37 vdd gnd cell_6t
Xbit_r38_c78 bl_78 br_78 wl_38 vdd gnd cell_6t
Xbit_r39_c78 bl_78 br_78 wl_39 vdd gnd cell_6t
Xbit_r40_c78 bl_78 br_78 wl_40 vdd gnd cell_6t
Xbit_r41_c78 bl_78 br_78 wl_41 vdd gnd cell_6t
Xbit_r42_c78 bl_78 br_78 wl_42 vdd gnd cell_6t
Xbit_r43_c78 bl_78 br_78 wl_43 vdd gnd cell_6t
Xbit_r44_c78 bl_78 br_78 wl_44 vdd gnd cell_6t
Xbit_r45_c78 bl_78 br_78 wl_45 vdd gnd cell_6t
Xbit_r46_c78 bl_78 br_78 wl_46 vdd gnd cell_6t
Xbit_r47_c78 bl_78 br_78 wl_47 vdd gnd cell_6t
Xbit_r48_c78 bl_78 br_78 wl_48 vdd gnd cell_6t
Xbit_r49_c78 bl_78 br_78 wl_49 vdd gnd cell_6t
Xbit_r50_c78 bl_78 br_78 wl_50 vdd gnd cell_6t
Xbit_r51_c78 bl_78 br_78 wl_51 vdd gnd cell_6t
Xbit_r52_c78 bl_78 br_78 wl_52 vdd gnd cell_6t
Xbit_r53_c78 bl_78 br_78 wl_53 vdd gnd cell_6t
Xbit_r54_c78 bl_78 br_78 wl_54 vdd gnd cell_6t
Xbit_r55_c78 bl_78 br_78 wl_55 vdd gnd cell_6t
Xbit_r56_c78 bl_78 br_78 wl_56 vdd gnd cell_6t
Xbit_r57_c78 bl_78 br_78 wl_57 vdd gnd cell_6t
Xbit_r58_c78 bl_78 br_78 wl_58 vdd gnd cell_6t
Xbit_r59_c78 bl_78 br_78 wl_59 vdd gnd cell_6t
Xbit_r60_c78 bl_78 br_78 wl_60 vdd gnd cell_6t
Xbit_r61_c78 bl_78 br_78 wl_61 vdd gnd cell_6t
Xbit_r62_c78 bl_78 br_78 wl_62 vdd gnd cell_6t
Xbit_r63_c78 bl_78 br_78 wl_63 vdd gnd cell_6t
Xbit_r64_c78 bl_78 br_78 wl_64 vdd gnd cell_6t
Xbit_r65_c78 bl_78 br_78 wl_65 vdd gnd cell_6t
Xbit_r66_c78 bl_78 br_78 wl_66 vdd gnd cell_6t
Xbit_r67_c78 bl_78 br_78 wl_67 vdd gnd cell_6t
Xbit_r68_c78 bl_78 br_78 wl_68 vdd gnd cell_6t
Xbit_r69_c78 bl_78 br_78 wl_69 vdd gnd cell_6t
Xbit_r70_c78 bl_78 br_78 wl_70 vdd gnd cell_6t
Xbit_r71_c78 bl_78 br_78 wl_71 vdd gnd cell_6t
Xbit_r72_c78 bl_78 br_78 wl_72 vdd gnd cell_6t
Xbit_r73_c78 bl_78 br_78 wl_73 vdd gnd cell_6t
Xbit_r74_c78 bl_78 br_78 wl_74 vdd gnd cell_6t
Xbit_r75_c78 bl_78 br_78 wl_75 vdd gnd cell_6t
Xbit_r76_c78 bl_78 br_78 wl_76 vdd gnd cell_6t
Xbit_r77_c78 bl_78 br_78 wl_77 vdd gnd cell_6t
Xbit_r78_c78 bl_78 br_78 wl_78 vdd gnd cell_6t
Xbit_r79_c78 bl_78 br_78 wl_79 vdd gnd cell_6t
Xbit_r80_c78 bl_78 br_78 wl_80 vdd gnd cell_6t
Xbit_r81_c78 bl_78 br_78 wl_81 vdd gnd cell_6t
Xbit_r82_c78 bl_78 br_78 wl_82 vdd gnd cell_6t
Xbit_r83_c78 bl_78 br_78 wl_83 vdd gnd cell_6t
Xbit_r84_c78 bl_78 br_78 wl_84 vdd gnd cell_6t
Xbit_r85_c78 bl_78 br_78 wl_85 vdd gnd cell_6t
Xbit_r86_c78 bl_78 br_78 wl_86 vdd gnd cell_6t
Xbit_r87_c78 bl_78 br_78 wl_87 vdd gnd cell_6t
Xbit_r88_c78 bl_78 br_78 wl_88 vdd gnd cell_6t
Xbit_r89_c78 bl_78 br_78 wl_89 vdd gnd cell_6t
Xbit_r90_c78 bl_78 br_78 wl_90 vdd gnd cell_6t
Xbit_r91_c78 bl_78 br_78 wl_91 vdd gnd cell_6t
Xbit_r92_c78 bl_78 br_78 wl_92 vdd gnd cell_6t
Xbit_r93_c78 bl_78 br_78 wl_93 vdd gnd cell_6t
Xbit_r94_c78 bl_78 br_78 wl_94 vdd gnd cell_6t
Xbit_r95_c78 bl_78 br_78 wl_95 vdd gnd cell_6t
Xbit_r96_c78 bl_78 br_78 wl_96 vdd gnd cell_6t
Xbit_r97_c78 bl_78 br_78 wl_97 vdd gnd cell_6t
Xbit_r98_c78 bl_78 br_78 wl_98 vdd gnd cell_6t
Xbit_r99_c78 bl_78 br_78 wl_99 vdd gnd cell_6t
Xbit_r100_c78 bl_78 br_78 wl_100 vdd gnd cell_6t
Xbit_r101_c78 bl_78 br_78 wl_101 vdd gnd cell_6t
Xbit_r102_c78 bl_78 br_78 wl_102 vdd gnd cell_6t
Xbit_r103_c78 bl_78 br_78 wl_103 vdd gnd cell_6t
Xbit_r104_c78 bl_78 br_78 wl_104 vdd gnd cell_6t
Xbit_r105_c78 bl_78 br_78 wl_105 vdd gnd cell_6t
Xbit_r106_c78 bl_78 br_78 wl_106 vdd gnd cell_6t
Xbit_r107_c78 bl_78 br_78 wl_107 vdd gnd cell_6t
Xbit_r108_c78 bl_78 br_78 wl_108 vdd gnd cell_6t
Xbit_r109_c78 bl_78 br_78 wl_109 vdd gnd cell_6t
Xbit_r110_c78 bl_78 br_78 wl_110 vdd gnd cell_6t
Xbit_r111_c78 bl_78 br_78 wl_111 vdd gnd cell_6t
Xbit_r112_c78 bl_78 br_78 wl_112 vdd gnd cell_6t
Xbit_r113_c78 bl_78 br_78 wl_113 vdd gnd cell_6t
Xbit_r114_c78 bl_78 br_78 wl_114 vdd gnd cell_6t
Xbit_r115_c78 bl_78 br_78 wl_115 vdd gnd cell_6t
Xbit_r116_c78 bl_78 br_78 wl_116 vdd gnd cell_6t
Xbit_r117_c78 bl_78 br_78 wl_117 vdd gnd cell_6t
Xbit_r118_c78 bl_78 br_78 wl_118 vdd gnd cell_6t
Xbit_r119_c78 bl_78 br_78 wl_119 vdd gnd cell_6t
Xbit_r120_c78 bl_78 br_78 wl_120 vdd gnd cell_6t
Xbit_r121_c78 bl_78 br_78 wl_121 vdd gnd cell_6t
Xbit_r122_c78 bl_78 br_78 wl_122 vdd gnd cell_6t
Xbit_r123_c78 bl_78 br_78 wl_123 vdd gnd cell_6t
Xbit_r124_c78 bl_78 br_78 wl_124 vdd gnd cell_6t
Xbit_r125_c78 bl_78 br_78 wl_125 vdd gnd cell_6t
Xbit_r126_c78 bl_78 br_78 wl_126 vdd gnd cell_6t
Xbit_r127_c78 bl_78 br_78 wl_127 vdd gnd cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd cell_6t
Xbit_r1_c79 bl_79 br_79 wl_1 vdd gnd cell_6t
Xbit_r2_c79 bl_79 br_79 wl_2 vdd gnd cell_6t
Xbit_r3_c79 bl_79 br_79 wl_3 vdd gnd cell_6t
Xbit_r4_c79 bl_79 br_79 wl_4 vdd gnd cell_6t
Xbit_r5_c79 bl_79 br_79 wl_5 vdd gnd cell_6t
Xbit_r6_c79 bl_79 br_79 wl_6 vdd gnd cell_6t
Xbit_r7_c79 bl_79 br_79 wl_7 vdd gnd cell_6t
Xbit_r8_c79 bl_79 br_79 wl_8 vdd gnd cell_6t
Xbit_r9_c79 bl_79 br_79 wl_9 vdd gnd cell_6t
Xbit_r10_c79 bl_79 br_79 wl_10 vdd gnd cell_6t
Xbit_r11_c79 bl_79 br_79 wl_11 vdd gnd cell_6t
Xbit_r12_c79 bl_79 br_79 wl_12 vdd gnd cell_6t
Xbit_r13_c79 bl_79 br_79 wl_13 vdd gnd cell_6t
Xbit_r14_c79 bl_79 br_79 wl_14 vdd gnd cell_6t
Xbit_r15_c79 bl_79 br_79 wl_15 vdd gnd cell_6t
Xbit_r16_c79 bl_79 br_79 wl_16 vdd gnd cell_6t
Xbit_r17_c79 bl_79 br_79 wl_17 vdd gnd cell_6t
Xbit_r18_c79 bl_79 br_79 wl_18 vdd gnd cell_6t
Xbit_r19_c79 bl_79 br_79 wl_19 vdd gnd cell_6t
Xbit_r20_c79 bl_79 br_79 wl_20 vdd gnd cell_6t
Xbit_r21_c79 bl_79 br_79 wl_21 vdd gnd cell_6t
Xbit_r22_c79 bl_79 br_79 wl_22 vdd gnd cell_6t
Xbit_r23_c79 bl_79 br_79 wl_23 vdd gnd cell_6t
Xbit_r24_c79 bl_79 br_79 wl_24 vdd gnd cell_6t
Xbit_r25_c79 bl_79 br_79 wl_25 vdd gnd cell_6t
Xbit_r26_c79 bl_79 br_79 wl_26 vdd gnd cell_6t
Xbit_r27_c79 bl_79 br_79 wl_27 vdd gnd cell_6t
Xbit_r28_c79 bl_79 br_79 wl_28 vdd gnd cell_6t
Xbit_r29_c79 bl_79 br_79 wl_29 vdd gnd cell_6t
Xbit_r30_c79 bl_79 br_79 wl_30 vdd gnd cell_6t
Xbit_r31_c79 bl_79 br_79 wl_31 vdd gnd cell_6t
Xbit_r32_c79 bl_79 br_79 wl_32 vdd gnd cell_6t
Xbit_r33_c79 bl_79 br_79 wl_33 vdd gnd cell_6t
Xbit_r34_c79 bl_79 br_79 wl_34 vdd gnd cell_6t
Xbit_r35_c79 bl_79 br_79 wl_35 vdd gnd cell_6t
Xbit_r36_c79 bl_79 br_79 wl_36 vdd gnd cell_6t
Xbit_r37_c79 bl_79 br_79 wl_37 vdd gnd cell_6t
Xbit_r38_c79 bl_79 br_79 wl_38 vdd gnd cell_6t
Xbit_r39_c79 bl_79 br_79 wl_39 vdd gnd cell_6t
Xbit_r40_c79 bl_79 br_79 wl_40 vdd gnd cell_6t
Xbit_r41_c79 bl_79 br_79 wl_41 vdd gnd cell_6t
Xbit_r42_c79 bl_79 br_79 wl_42 vdd gnd cell_6t
Xbit_r43_c79 bl_79 br_79 wl_43 vdd gnd cell_6t
Xbit_r44_c79 bl_79 br_79 wl_44 vdd gnd cell_6t
Xbit_r45_c79 bl_79 br_79 wl_45 vdd gnd cell_6t
Xbit_r46_c79 bl_79 br_79 wl_46 vdd gnd cell_6t
Xbit_r47_c79 bl_79 br_79 wl_47 vdd gnd cell_6t
Xbit_r48_c79 bl_79 br_79 wl_48 vdd gnd cell_6t
Xbit_r49_c79 bl_79 br_79 wl_49 vdd gnd cell_6t
Xbit_r50_c79 bl_79 br_79 wl_50 vdd gnd cell_6t
Xbit_r51_c79 bl_79 br_79 wl_51 vdd gnd cell_6t
Xbit_r52_c79 bl_79 br_79 wl_52 vdd gnd cell_6t
Xbit_r53_c79 bl_79 br_79 wl_53 vdd gnd cell_6t
Xbit_r54_c79 bl_79 br_79 wl_54 vdd gnd cell_6t
Xbit_r55_c79 bl_79 br_79 wl_55 vdd gnd cell_6t
Xbit_r56_c79 bl_79 br_79 wl_56 vdd gnd cell_6t
Xbit_r57_c79 bl_79 br_79 wl_57 vdd gnd cell_6t
Xbit_r58_c79 bl_79 br_79 wl_58 vdd gnd cell_6t
Xbit_r59_c79 bl_79 br_79 wl_59 vdd gnd cell_6t
Xbit_r60_c79 bl_79 br_79 wl_60 vdd gnd cell_6t
Xbit_r61_c79 bl_79 br_79 wl_61 vdd gnd cell_6t
Xbit_r62_c79 bl_79 br_79 wl_62 vdd gnd cell_6t
Xbit_r63_c79 bl_79 br_79 wl_63 vdd gnd cell_6t
Xbit_r64_c79 bl_79 br_79 wl_64 vdd gnd cell_6t
Xbit_r65_c79 bl_79 br_79 wl_65 vdd gnd cell_6t
Xbit_r66_c79 bl_79 br_79 wl_66 vdd gnd cell_6t
Xbit_r67_c79 bl_79 br_79 wl_67 vdd gnd cell_6t
Xbit_r68_c79 bl_79 br_79 wl_68 vdd gnd cell_6t
Xbit_r69_c79 bl_79 br_79 wl_69 vdd gnd cell_6t
Xbit_r70_c79 bl_79 br_79 wl_70 vdd gnd cell_6t
Xbit_r71_c79 bl_79 br_79 wl_71 vdd gnd cell_6t
Xbit_r72_c79 bl_79 br_79 wl_72 vdd gnd cell_6t
Xbit_r73_c79 bl_79 br_79 wl_73 vdd gnd cell_6t
Xbit_r74_c79 bl_79 br_79 wl_74 vdd gnd cell_6t
Xbit_r75_c79 bl_79 br_79 wl_75 vdd gnd cell_6t
Xbit_r76_c79 bl_79 br_79 wl_76 vdd gnd cell_6t
Xbit_r77_c79 bl_79 br_79 wl_77 vdd gnd cell_6t
Xbit_r78_c79 bl_79 br_79 wl_78 vdd gnd cell_6t
Xbit_r79_c79 bl_79 br_79 wl_79 vdd gnd cell_6t
Xbit_r80_c79 bl_79 br_79 wl_80 vdd gnd cell_6t
Xbit_r81_c79 bl_79 br_79 wl_81 vdd gnd cell_6t
Xbit_r82_c79 bl_79 br_79 wl_82 vdd gnd cell_6t
Xbit_r83_c79 bl_79 br_79 wl_83 vdd gnd cell_6t
Xbit_r84_c79 bl_79 br_79 wl_84 vdd gnd cell_6t
Xbit_r85_c79 bl_79 br_79 wl_85 vdd gnd cell_6t
Xbit_r86_c79 bl_79 br_79 wl_86 vdd gnd cell_6t
Xbit_r87_c79 bl_79 br_79 wl_87 vdd gnd cell_6t
Xbit_r88_c79 bl_79 br_79 wl_88 vdd gnd cell_6t
Xbit_r89_c79 bl_79 br_79 wl_89 vdd gnd cell_6t
Xbit_r90_c79 bl_79 br_79 wl_90 vdd gnd cell_6t
Xbit_r91_c79 bl_79 br_79 wl_91 vdd gnd cell_6t
Xbit_r92_c79 bl_79 br_79 wl_92 vdd gnd cell_6t
Xbit_r93_c79 bl_79 br_79 wl_93 vdd gnd cell_6t
Xbit_r94_c79 bl_79 br_79 wl_94 vdd gnd cell_6t
Xbit_r95_c79 bl_79 br_79 wl_95 vdd gnd cell_6t
Xbit_r96_c79 bl_79 br_79 wl_96 vdd gnd cell_6t
Xbit_r97_c79 bl_79 br_79 wl_97 vdd gnd cell_6t
Xbit_r98_c79 bl_79 br_79 wl_98 vdd gnd cell_6t
Xbit_r99_c79 bl_79 br_79 wl_99 vdd gnd cell_6t
Xbit_r100_c79 bl_79 br_79 wl_100 vdd gnd cell_6t
Xbit_r101_c79 bl_79 br_79 wl_101 vdd gnd cell_6t
Xbit_r102_c79 bl_79 br_79 wl_102 vdd gnd cell_6t
Xbit_r103_c79 bl_79 br_79 wl_103 vdd gnd cell_6t
Xbit_r104_c79 bl_79 br_79 wl_104 vdd gnd cell_6t
Xbit_r105_c79 bl_79 br_79 wl_105 vdd gnd cell_6t
Xbit_r106_c79 bl_79 br_79 wl_106 vdd gnd cell_6t
Xbit_r107_c79 bl_79 br_79 wl_107 vdd gnd cell_6t
Xbit_r108_c79 bl_79 br_79 wl_108 vdd gnd cell_6t
Xbit_r109_c79 bl_79 br_79 wl_109 vdd gnd cell_6t
Xbit_r110_c79 bl_79 br_79 wl_110 vdd gnd cell_6t
Xbit_r111_c79 bl_79 br_79 wl_111 vdd gnd cell_6t
Xbit_r112_c79 bl_79 br_79 wl_112 vdd gnd cell_6t
Xbit_r113_c79 bl_79 br_79 wl_113 vdd gnd cell_6t
Xbit_r114_c79 bl_79 br_79 wl_114 vdd gnd cell_6t
Xbit_r115_c79 bl_79 br_79 wl_115 vdd gnd cell_6t
Xbit_r116_c79 bl_79 br_79 wl_116 vdd gnd cell_6t
Xbit_r117_c79 bl_79 br_79 wl_117 vdd gnd cell_6t
Xbit_r118_c79 bl_79 br_79 wl_118 vdd gnd cell_6t
Xbit_r119_c79 bl_79 br_79 wl_119 vdd gnd cell_6t
Xbit_r120_c79 bl_79 br_79 wl_120 vdd gnd cell_6t
Xbit_r121_c79 bl_79 br_79 wl_121 vdd gnd cell_6t
Xbit_r122_c79 bl_79 br_79 wl_122 vdd gnd cell_6t
Xbit_r123_c79 bl_79 br_79 wl_123 vdd gnd cell_6t
Xbit_r124_c79 bl_79 br_79 wl_124 vdd gnd cell_6t
Xbit_r125_c79 bl_79 br_79 wl_125 vdd gnd cell_6t
Xbit_r126_c79 bl_79 br_79 wl_126 vdd gnd cell_6t
Xbit_r127_c79 bl_79 br_79 wl_127 vdd gnd cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd cell_6t
Xbit_r1_c80 bl_80 br_80 wl_1 vdd gnd cell_6t
Xbit_r2_c80 bl_80 br_80 wl_2 vdd gnd cell_6t
Xbit_r3_c80 bl_80 br_80 wl_3 vdd gnd cell_6t
Xbit_r4_c80 bl_80 br_80 wl_4 vdd gnd cell_6t
Xbit_r5_c80 bl_80 br_80 wl_5 vdd gnd cell_6t
Xbit_r6_c80 bl_80 br_80 wl_6 vdd gnd cell_6t
Xbit_r7_c80 bl_80 br_80 wl_7 vdd gnd cell_6t
Xbit_r8_c80 bl_80 br_80 wl_8 vdd gnd cell_6t
Xbit_r9_c80 bl_80 br_80 wl_9 vdd gnd cell_6t
Xbit_r10_c80 bl_80 br_80 wl_10 vdd gnd cell_6t
Xbit_r11_c80 bl_80 br_80 wl_11 vdd gnd cell_6t
Xbit_r12_c80 bl_80 br_80 wl_12 vdd gnd cell_6t
Xbit_r13_c80 bl_80 br_80 wl_13 vdd gnd cell_6t
Xbit_r14_c80 bl_80 br_80 wl_14 vdd gnd cell_6t
Xbit_r15_c80 bl_80 br_80 wl_15 vdd gnd cell_6t
Xbit_r16_c80 bl_80 br_80 wl_16 vdd gnd cell_6t
Xbit_r17_c80 bl_80 br_80 wl_17 vdd gnd cell_6t
Xbit_r18_c80 bl_80 br_80 wl_18 vdd gnd cell_6t
Xbit_r19_c80 bl_80 br_80 wl_19 vdd gnd cell_6t
Xbit_r20_c80 bl_80 br_80 wl_20 vdd gnd cell_6t
Xbit_r21_c80 bl_80 br_80 wl_21 vdd gnd cell_6t
Xbit_r22_c80 bl_80 br_80 wl_22 vdd gnd cell_6t
Xbit_r23_c80 bl_80 br_80 wl_23 vdd gnd cell_6t
Xbit_r24_c80 bl_80 br_80 wl_24 vdd gnd cell_6t
Xbit_r25_c80 bl_80 br_80 wl_25 vdd gnd cell_6t
Xbit_r26_c80 bl_80 br_80 wl_26 vdd gnd cell_6t
Xbit_r27_c80 bl_80 br_80 wl_27 vdd gnd cell_6t
Xbit_r28_c80 bl_80 br_80 wl_28 vdd gnd cell_6t
Xbit_r29_c80 bl_80 br_80 wl_29 vdd gnd cell_6t
Xbit_r30_c80 bl_80 br_80 wl_30 vdd gnd cell_6t
Xbit_r31_c80 bl_80 br_80 wl_31 vdd gnd cell_6t
Xbit_r32_c80 bl_80 br_80 wl_32 vdd gnd cell_6t
Xbit_r33_c80 bl_80 br_80 wl_33 vdd gnd cell_6t
Xbit_r34_c80 bl_80 br_80 wl_34 vdd gnd cell_6t
Xbit_r35_c80 bl_80 br_80 wl_35 vdd gnd cell_6t
Xbit_r36_c80 bl_80 br_80 wl_36 vdd gnd cell_6t
Xbit_r37_c80 bl_80 br_80 wl_37 vdd gnd cell_6t
Xbit_r38_c80 bl_80 br_80 wl_38 vdd gnd cell_6t
Xbit_r39_c80 bl_80 br_80 wl_39 vdd gnd cell_6t
Xbit_r40_c80 bl_80 br_80 wl_40 vdd gnd cell_6t
Xbit_r41_c80 bl_80 br_80 wl_41 vdd gnd cell_6t
Xbit_r42_c80 bl_80 br_80 wl_42 vdd gnd cell_6t
Xbit_r43_c80 bl_80 br_80 wl_43 vdd gnd cell_6t
Xbit_r44_c80 bl_80 br_80 wl_44 vdd gnd cell_6t
Xbit_r45_c80 bl_80 br_80 wl_45 vdd gnd cell_6t
Xbit_r46_c80 bl_80 br_80 wl_46 vdd gnd cell_6t
Xbit_r47_c80 bl_80 br_80 wl_47 vdd gnd cell_6t
Xbit_r48_c80 bl_80 br_80 wl_48 vdd gnd cell_6t
Xbit_r49_c80 bl_80 br_80 wl_49 vdd gnd cell_6t
Xbit_r50_c80 bl_80 br_80 wl_50 vdd gnd cell_6t
Xbit_r51_c80 bl_80 br_80 wl_51 vdd gnd cell_6t
Xbit_r52_c80 bl_80 br_80 wl_52 vdd gnd cell_6t
Xbit_r53_c80 bl_80 br_80 wl_53 vdd gnd cell_6t
Xbit_r54_c80 bl_80 br_80 wl_54 vdd gnd cell_6t
Xbit_r55_c80 bl_80 br_80 wl_55 vdd gnd cell_6t
Xbit_r56_c80 bl_80 br_80 wl_56 vdd gnd cell_6t
Xbit_r57_c80 bl_80 br_80 wl_57 vdd gnd cell_6t
Xbit_r58_c80 bl_80 br_80 wl_58 vdd gnd cell_6t
Xbit_r59_c80 bl_80 br_80 wl_59 vdd gnd cell_6t
Xbit_r60_c80 bl_80 br_80 wl_60 vdd gnd cell_6t
Xbit_r61_c80 bl_80 br_80 wl_61 vdd gnd cell_6t
Xbit_r62_c80 bl_80 br_80 wl_62 vdd gnd cell_6t
Xbit_r63_c80 bl_80 br_80 wl_63 vdd gnd cell_6t
Xbit_r64_c80 bl_80 br_80 wl_64 vdd gnd cell_6t
Xbit_r65_c80 bl_80 br_80 wl_65 vdd gnd cell_6t
Xbit_r66_c80 bl_80 br_80 wl_66 vdd gnd cell_6t
Xbit_r67_c80 bl_80 br_80 wl_67 vdd gnd cell_6t
Xbit_r68_c80 bl_80 br_80 wl_68 vdd gnd cell_6t
Xbit_r69_c80 bl_80 br_80 wl_69 vdd gnd cell_6t
Xbit_r70_c80 bl_80 br_80 wl_70 vdd gnd cell_6t
Xbit_r71_c80 bl_80 br_80 wl_71 vdd gnd cell_6t
Xbit_r72_c80 bl_80 br_80 wl_72 vdd gnd cell_6t
Xbit_r73_c80 bl_80 br_80 wl_73 vdd gnd cell_6t
Xbit_r74_c80 bl_80 br_80 wl_74 vdd gnd cell_6t
Xbit_r75_c80 bl_80 br_80 wl_75 vdd gnd cell_6t
Xbit_r76_c80 bl_80 br_80 wl_76 vdd gnd cell_6t
Xbit_r77_c80 bl_80 br_80 wl_77 vdd gnd cell_6t
Xbit_r78_c80 bl_80 br_80 wl_78 vdd gnd cell_6t
Xbit_r79_c80 bl_80 br_80 wl_79 vdd gnd cell_6t
Xbit_r80_c80 bl_80 br_80 wl_80 vdd gnd cell_6t
Xbit_r81_c80 bl_80 br_80 wl_81 vdd gnd cell_6t
Xbit_r82_c80 bl_80 br_80 wl_82 vdd gnd cell_6t
Xbit_r83_c80 bl_80 br_80 wl_83 vdd gnd cell_6t
Xbit_r84_c80 bl_80 br_80 wl_84 vdd gnd cell_6t
Xbit_r85_c80 bl_80 br_80 wl_85 vdd gnd cell_6t
Xbit_r86_c80 bl_80 br_80 wl_86 vdd gnd cell_6t
Xbit_r87_c80 bl_80 br_80 wl_87 vdd gnd cell_6t
Xbit_r88_c80 bl_80 br_80 wl_88 vdd gnd cell_6t
Xbit_r89_c80 bl_80 br_80 wl_89 vdd gnd cell_6t
Xbit_r90_c80 bl_80 br_80 wl_90 vdd gnd cell_6t
Xbit_r91_c80 bl_80 br_80 wl_91 vdd gnd cell_6t
Xbit_r92_c80 bl_80 br_80 wl_92 vdd gnd cell_6t
Xbit_r93_c80 bl_80 br_80 wl_93 vdd gnd cell_6t
Xbit_r94_c80 bl_80 br_80 wl_94 vdd gnd cell_6t
Xbit_r95_c80 bl_80 br_80 wl_95 vdd gnd cell_6t
Xbit_r96_c80 bl_80 br_80 wl_96 vdd gnd cell_6t
Xbit_r97_c80 bl_80 br_80 wl_97 vdd gnd cell_6t
Xbit_r98_c80 bl_80 br_80 wl_98 vdd gnd cell_6t
Xbit_r99_c80 bl_80 br_80 wl_99 vdd gnd cell_6t
Xbit_r100_c80 bl_80 br_80 wl_100 vdd gnd cell_6t
Xbit_r101_c80 bl_80 br_80 wl_101 vdd gnd cell_6t
Xbit_r102_c80 bl_80 br_80 wl_102 vdd gnd cell_6t
Xbit_r103_c80 bl_80 br_80 wl_103 vdd gnd cell_6t
Xbit_r104_c80 bl_80 br_80 wl_104 vdd gnd cell_6t
Xbit_r105_c80 bl_80 br_80 wl_105 vdd gnd cell_6t
Xbit_r106_c80 bl_80 br_80 wl_106 vdd gnd cell_6t
Xbit_r107_c80 bl_80 br_80 wl_107 vdd gnd cell_6t
Xbit_r108_c80 bl_80 br_80 wl_108 vdd gnd cell_6t
Xbit_r109_c80 bl_80 br_80 wl_109 vdd gnd cell_6t
Xbit_r110_c80 bl_80 br_80 wl_110 vdd gnd cell_6t
Xbit_r111_c80 bl_80 br_80 wl_111 vdd gnd cell_6t
Xbit_r112_c80 bl_80 br_80 wl_112 vdd gnd cell_6t
Xbit_r113_c80 bl_80 br_80 wl_113 vdd gnd cell_6t
Xbit_r114_c80 bl_80 br_80 wl_114 vdd gnd cell_6t
Xbit_r115_c80 bl_80 br_80 wl_115 vdd gnd cell_6t
Xbit_r116_c80 bl_80 br_80 wl_116 vdd gnd cell_6t
Xbit_r117_c80 bl_80 br_80 wl_117 vdd gnd cell_6t
Xbit_r118_c80 bl_80 br_80 wl_118 vdd gnd cell_6t
Xbit_r119_c80 bl_80 br_80 wl_119 vdd gnd cell_6t
Xbit_r120_c80 bl_80 br_80 wl_120 vdd gnd cell_6t
Xbit_r121_c80 bl_80 br_80 wl_121 vdd gnd cell_6t
Xbit_r122_c80 bl_80 br_80 wl_122 vdd gnd cell_6t
Xbit_r123_c80 bl_80 br_80 wl_123 vdd gnd cell_6t
Xbit_r124_c80 bl_80 br_80 wl_124 vdd gnd cell_6t
Xbit_r125_c80 bl_80 br_80 wl_125 vdd gnd cell_6t
Xbit_r126_c80 bl_80 br_80 wl_126 vdd gnd cell_6t
Xbit_r127_c80 bl_80 br_80 wl_127 vdd gnd cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd cell_6t
Xbit_r1_c81 bl_81 br_81 wl_1 vdd gnd cell_6t
Xbit_r2_c81 bl_81 br_81 wl_2 vdd gnd cell_6t
Xbit_r3_c81 bl_81 br_81 wl_3 vdd gnd cell_6t
Xbit_r4_c81 bl_81 br_81 wl_4 vdd gnd cell_6t
Xbit_r5_c81 bl_81 br_81 wl_5 vdd gnd cell_6t
Xbit_r6_c81 bl_81 br_81 wl_6 vdd gnd cell_6t
Xbit_r7_c81 bl_81 br_81 wl_7 vdd gnd cell_6t
Xbit_r8_c81 bl_81 br_81 wl_8 vdd gnd cell_6t
Xbit_r9_c81 bl_81 br_81 wl_9 vdd gnd cell_6t
Xbit_r10_c81 bl_81 br_81 wl_10 vdd gnd cell_6t
Xbit_r11_c81 bl_81 br_81 wl_11 vdd gnd cell_6t
Xbit_r12_c81 bl_81 br_81 wl_12 vdd gnd cell_6t
Xbit_r13_c81 bl_81 br_81 wl_13 vdd gnd cell_6t
Xbit_r14_c81 bl_81 br_81 wl_14 vdd gnd cell_6t
Xbit_r15_c81 bl_81 br_81 wl_15 vdd gnd cell_6t
Xbit_r16_c81 bl_81 br_81 wl_16 vdd gnd cell_6t
Xbit_r17_c81 bl_81 br_81 wl_17 vdd gnd cell_6t
Xbit_r18_c81 bl_81 br_81 wl_18 vdd gnd cell_6t
Xbit_r19_c81 bl_81 br_81 wl_19 vdd gnd cell_6t
Xbit_r20_c81 bl_81 br_81 wl_20 vdd gnd cell_6t
Xbit_r21_c81 bl_81 br_81 wl_21 vdd gnd cell_6t
Xbit_r22_c81 bl_81 br_81 wl_22 vdd gnd cell_6t
Xbit_r23_c81 bl_81 br_81 wl_23 vdd gnd cell_6t
Xbit_r24_c81 bl_81 br_81 wl_24 vdd gnd cell_6t
Xbit_r25_c81 bl_81 br_81 wl_25 vdd gnd cell_6t
Xbit_r26_c81 bl_81 br_81 wl_26 vdd gnd cell_6t
Xbit_r27_c81 bl_81 br_81 wl_27 vdd gnd cell_6t
Xbit_r28_c81 bl_81 br_81 wl_28 vdd gnd cell_6t
Xbit_r29_c81 bl_81 br_81 wl_29 vdd gnd cell_6t
Xbit_r30_c81 bl_81 br_81 wl_30 vdd gnd cell_6t
Xbit_r31_c81 bl_81 br_81 wl_31 vdd gnd cell_6t
Xbit_r32_c81 bl_81 br_81 wl_32 vdd gnd cell_6t
Xbit_r33_c81 bl_81 br_81 wl_33 vdd gnd cell_6t
Xbit_r34_c81 bl_81 br_81 wl_34 vdd gnd cell_6t
Xbit_r35_c81 bl_81 br_81 wl_35 vdd gnd cell_6t
Xbit_r36_c81 bl_81 br_81 wl_36 vdd gnd cell_6t
Xbit_r37_c81 bl_81 br_81 wl_37 vdd gnd cell_6t
Xbit_r38_c81 bl_81 br_81 wl_38 vdd gnd cell_6t
Xbit_r39_c81 bl_81 br_81 wl_39 vdd gnd cell_6t
Xbit_r40_c81 bl_81 br_81 wl_40 vdd gnd cell_6t
Xbit_r41_c81 bl_81 br_81 wl_41 vdd gnd cell_6t
Xbit_r42_c81 bl_81 br_81 wl_42 vdd gnd cell_6t
Xbit_r43_c81 bl_81 br_81 wl_43 vdd gnd cell_6t
Xbit_r44_c81 bl_81 br_81 wl_44 vdd gnd cell_6t
Xbit_r45_c81 bl_81 br_81 wl_45 vdd gnd cell_6t
Xbit_r46_c81 bl_81 br_81 wl_46 vdd gnd cell_6t
Xbit_r47_c81 bl_81 br_81 wl_47 vdd gnd cell_6t
Xbit_r48_c81 bl_81 br_81 wl_48 vdd gnd cell_6t
Xbit_r49_c81 bl_81 br_81 wl_49 vdd gnd cell_6t
Xbit_r50_c81 bl_81 br_81 wl_50 vdd gnd cell_6t
Xbit_r51_c81 bl_81 br_81 wl_51 vdd gnd cell_6t
Xbit_r52_c81 bl_81 br_81 wl_52 vdd gnd cell_6t
Xbit_r53_c81 bl_81 br_81 wl_53 vdd gnd cell_6t
Xbit_r54_c81 bl_81 br_81 wl_54 vdd gnd cell_6t
Xbit_r55_c81 bl_81 br_81 wl_55 vdd gnd cell_6t
Xbit_r56_c81 bl_81 br_81 wl_56 vdd gnd cell_6t
Xbit_r57_c81 bl_81 br_81 wl_57 vdd gnd cell_6t
Xbit_r58_c81 bl_81 br_81 wl_58 vdd gnd cell_6t
Xbit_r59_c81 bl_81 br_81 wl_59 vdd gnd cell_6t
Xbit_r60_c81 bl_81 br_81 wl_60 vdd gnd cell_6t
Xbit_r61_c81 bl_81 br_81 wl_61 vdd gnd cell_6t
Xbit_r62_c81 bl_81 br_81 wl_62 vdd gnd cell_6t
Xbit_r63_c81 bl_81 br_81 wl_63 vdd gnd cell_6t
Xbit_r64_c81 bl_81 br_81 wl_64 vdd gnd cell_6t
Xbit_r65_c81 bl_81 br_81 wl_65 vdd gnd cell_6t
Xbit_r66_c81 bl_81 br_81 wl_66 vdd gnd cell_6t
Xbit_r67_c81 bl_81 br_81 wl_67 vdd gnd cell_6t
Xbit_r68_c81 bl_81 br_81 wl_68 vdd gnd cell_6t
Xbit_r69_c81 bl_81 br_81 wl_69 vdd gnd cell_6t
Xbit_r70_c81 bl_81 br_81 wl_70 vdd gnd cell_6t
Xbit_r71_c81 bl_81 br_81 wl_71 vdd gnd cell_6t
Xbit_r72_c81 bl_81 br_81 wl_72 vdd gnd cell_6t
Xbit_r73_c81 bl_81 br_81 wl_73 vdd gnd cell_6t
Xbit_r74_c81 bl_81 br_81 wl_74 vdd gnd cell_6t
Xbit_r75_c81 bl_81 br_81 wl_75 vdd gnd cell_6t
Xbit_r76_c81 bl_81 br_81 wl_76 vdd gnd cell_6t
Xbit_r77_c81 bl_81 br_81 wl_77 vdd gnd cell_6t
Xbit_r78_c81 bl_81 br_81 wl_78 vdd gnd cell_6t
Xbit_r79_c81 bl_81 br_81 wl_79 vdd gnd cell_6t
Xbit_r80_c81 bl_81 br_81 wl_80 vdd gnd cell_6t
Xbit_r81_c81 bl_81 br_81 wl_81 vdd gnd cell_6t
Xbit_r82_c81 bl_81 br_81 wl_82 vdd gnd cell_6t
Xbit_r83_c81 bl_81 br_81 wl_83 vdd gnd cell_6t
Xbit_r84_c81 bl_81 br_81 wl_84 vdd gnd cell_6t
Xbit_r85_c81 bl_81 br_81 wl_85 vdd gnd cell_6t
Xbit_r86_c81 bl_81 br_81 wl_86 vdd gnd cell_6t
Xbit_r87_c81 bl_81 br_81 wl_87 vdd gnd cell_6t
Xbit_r88_c81 bl_81 br_81 wl_88 vdd gnd cell_6t
Xbit_r89_c81 bl_81 br_81 wl_89 vdd gnd cell_6t
Xbit_r90_c81 bl_81 br_81 wl_90 vdd gnd cell_6t
Xbit_r91_c81 bl_81 br_81 wl_91 vdd gnd cell_6t
Xbit_r92_c81 bl_81 br_81 wl_92 vdd gnd cell_6t
Xbit_r93_c81 bl_81 br_81 wl_93 vdd gnd cell_6t
Xbit_r94_c81 bl_81 br_81 wl_94 vdd gnd cell_6t
Xbit_r95_c81 bl_81 br_81 wl_95 vdd gnd cell_6t
Xbit_r96_c81 bl_81 br_81 wl_96 vdd gnd cell_6t
Xbit_r97_c81 bl_81 br_81 wl_97 vdd gnd cell_6t
Xbit_r98_c81 bl_81 br_81 wl_98 vdd gnd cell_6t
Xbit_r99_c81 bl_81 br_81 wl_99 vdd gnd cell_6t
Xbit_r100_c81 bl_81 br_81 wl_100 vdd gnd cell_6t
Xbit_r101_c81 bl_81 br_81 wl_101 vdd gnd cell_6t
Xbit_r102_c81 bl_81 br_81 wl_102 vdd gnd cell_6t
Xbit_r103_c81 bl_81 br_81 wl_103 vdd gnd cell_6t
Xbit_r104_c81 bl_81 br_81 wl_104 vdd gnd cell_6t
Xbit_r105_c81 bl_81 br_81 wl_105 vdd gnd cell_6t
Xbit_r106_c81 bl_81 br_81 wl_106 vdd gnd cell_6t
Xbit_r107_c81 bl_81 br_81 wl_107 vdd gnd cell_6t
Xbit_r108_c81 bl_81 br_81 wl_108 vdd gnd cell_6t
Xbit_r109_c81 bl_81 br_81 wl_109 vdd gnd cell_6t
Xbit_r110_c81 bl_81 br_81 wl_110 vdd gnd cell_6t
Xbit_r111_c81 bl_81 br_81 wl_111 vdd gnd cell_6t
Xbit_r112_c81 bl_81 br_81 wl_112 vdd gnd cell_6t
Xbit_r113_c81 bl_81 br_81 wl_113 vdd gnd cell_6t
Xbit_r114_c81 bl_81 br_81 wl_114 vdd gnd cell_6t
Xbit_r115_c81 bl_81 br_81 wl_115 vdd gnd cell_6t
Xbit_r116_c81 bl_81 br_81 wl_116 vdd gnd cell_6t
Xbit_r117_c81 bl_81 br_81 wl_117 vdd gnd cell_6t
Xbit_r118_c81 bl_81 br_81 wl_118 vdd gnd cell_6t
Xbit_r119_c81 bl_81 br_81 wl_119 vdd gnd cell_6t
Xbit_r120_c81 bl_81 br_81 wl_120 vdd gnd cell_6t
Xbit_r121_c81 bl_81 br_81 wl_121 vdd gnd cell_6t
Xbit_r122_c81 bl_81 br_81 wl_122 vdd gnd cell_6t
Xbit_r123_c81 bl_81 br_81 wl_123 vdd gnd cell_6t
Xbit_r124_c81 bl_81 br_81 wl_124 vdd gnd cell_6t
Xbit_r125_c81 bl_81 br_81 wl_125 vdd gnd cell_6t
Xbit_r126_c81 bl_81 br_81 wl_126 vdd gnd cell_6t
Xbit_r127_c81 bl_81 br_81 wl_127 vdd gnd cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd cell_6t
Xbit_r1_c82 bl_82 br_82 wl_1 vdd gnd cell_6t
Xbit_r2_c82 bl_82 br_82 wl_2 vdd gnd cell_6t
Xbit_r3_c82 bl_82 br_82 wl_3 vdd gnd cell_6t
Xbit_r4_c82 bl_82 br_82 wl_4 vdd gnd cell_6t
Xbit_r5_c82 bl_82 br_82 wl_5 vdd gnd cell_6t
Xbit_r6_c82 bl_82 br_82 wl_6 vdd gnd cell_6t
Xbit_r7_c82 bl_82 br_82 wl_7 vdd gnd cell_6t
Xbit_r8_c82 bl_82 br_82 wl_8 vdd gnd cell_6t
Xbit_r9_c82 bl_82 br_82 wl_9 vdd gnd cell_6t
Xbit_r10_c82 bl_82 br_82 wl_10 vdd gnd cell_6t
Xbit_r11_c82 bl_82 br_82 wl_11 vdd gnd cell_6t
Xbit_r12_c82 bl_82 br_82 wl_12 vdd gnd cell_6t
Xbit_r13_c82 bl_82 br_82 wl_13 vdd gnd cell_6t
Xbit_r14_c82 bl_82 br_82 wl_14 vdd gnd cell_6t
Xbit_r15_c82 bl_82 br_82 wl_15 vdd gnd cell_6t
Xbit_r16_c82 bl_82 br_82 wl_16 vdd gnd cell_6t
Xbit_r17_c82 bl_82 br_82 wl_17 vdd gnd cell_6t
Xbit_r18_c82 bl_82 br_82 wl_18 vdd gnd cell_6t
Xbit_r19_c82 bl_82 br_82 wl_19 vdd gnd cell_6t
Xbit_r20_c82 bl_82 br_82 wl_20 vdd gnd cell_6t
Xbit_r21_c82 bl_82 br_82 wl_21 vdd gnd cell_6t
Xbit_r22_c82 bl_82 br_82 wl_22 vdd gnd cell_6t
Xbit_r23_c82 bl_82 br_82 wl_23 vdd gnd cell_6t
Xbit_r24_c82 bl_82 br_82 wl_24 vdd gnd cell_6t
Xbit_r25_c82 bl_82 br_82 wl_25 vdd gnd cell_6t
Xbit_r26_c82 bl_82 br_82 wl_26 vdd gnd cell_6t
Xbit_r27_c82 bl_82 br_82 wl_27 vdd gnd cell_6t
Xbit_r28_c82 bl_82 br_82 wl_28 vdd gnd cell_6t
Xbit_r29_c82 bl_82 br_82 wl_29 vdd gnd cell_6t
Xbit_r30_c82 bl_82 br_82 wl_30 vdd gnd cell_6t
Xbit_r31_c82 bl_82 br_82 wl_31 vdd gnd cell_6t
Xbit_r32_c82 bl_82 br_82 wl_32 vdd gnd cell_6t
Xbit_r33_c82 bl_82 br_82 wl_33 vdd gnd cell_6t
Xbit_r34_c82 bl_82 br_82 wl_34 vdd gnd cell_6t
Xbit_r35_c82 bl_82 br_82 wl_35 vdd gnd cell_6t
Xbit_r36_c82 bl_82 br_82 wl_36 vdd gnd cell_6t
Xbit_r37_c82 bl_82 br_82 wl_37 vdd gnd cell_6t
Xbit_r38_c82 bl_82 br_82 wl_38 vdd gnd cell_6t
Xbit_r39_c82 bl_82 br_82 wl_39 vdd gnd cell_6t
Xbit_r40_c82 bl_82 br_82 wl_40 vdd gnd cell_6t
Xbit_r41_c82 bl_82 br_82 wl_41 vdd gnd cell_6t
Xbit_r42_c82 bl_82 br_82 wl_42 vdd gnd cell_6t
Xbit_r43_c82 bl_82 br_82 wl_43 vdd gnd cell_6t
Xbit_r44_c82 bl_82 br_82 wl_44 vdd gnd cell_6t
Xbit_r45_c82 bl_82 br_82 wl_45 vdd gnd cell_6t
Xbit_r46_c82 bl_82 br_82 wl_46 vdd gnd cell_6t
Xbit_r47_c82 bl_82 br_82 wl_47 vdd gnd cell_6t
Xbit_r48_c82 bl_82 br_82 wl_48 vdd gnd cell_6t
Xbit_r49_c82 bl_82 br_82 wl_49 vdd gnd cell_6t
Xbit_r50_c82 bl_82 br_82 wl_50 vdd gnd cell_6t
Xbit_r51_c82 bl_82 br_82 wl_51 vdd gnd cell_6t
Xbit_r52_c82 bl_82 br_82 wl_52 vdd gnd cell_6t
Xbit_r53_c82 bl_82 br_82 wl_53 vdd gnd cell_6t
Xbit_r54_c82 bl_82 br_82 wl_54 vdd gnd cell_6t
Xbit_r55_c82 bl_82 br_82 wl_55 vdd gnd cell_6t
Xbit_r56_c82 bl_82 br_82 wl_56 vdd gnd cell_6t
Xbit_r57_c82 bl_82 br_82 wl_57 vdd gnd cell_6t
Xbit_r58_c82 bl_82 br_82 wl_58 vdd gnd cell_6t
Xbit_r59_c82 bl_82 br_82 wl_59 vdd gnd cell_6t
Xbit_r60_c82 bl_82 br_82 wl_60 vdd gnd cell_6t
Xbit_r61_c82 bl_82 br_82 wl_61 vdd gnd cell_6t
Xbit_r62_c82 bl_82 br_82 wl_62 vdd gnd cell_6t
Xbit_r63_c82 bl_82 br_82 wl_63 vdd gnd cell_6t
Xbit_r64_c82 bl_82 br_82 wl_64 vdd gnd cell_6t
Xbit_r65_c82 bl_82 br_82 wl_65 vdd gnd cell_6t
Xbit_r66_c82 bl_82 br_82 wl_66 vdd gnd cell_6t
Xbit_r67_c82 bl_82 br_82 wl_67 vdd gnd cell_6t
Xbit_r68_c82 bl_82 br_82 wl_68 vdd gnd cell_6t
Xbit_r69_c82 bl_82 br_82 wl_69 vdd gnd cell_6t
Xbit_r70_c82 bl_82 br_82 wl_70 vdd gnd cell_6t
Xbit_r71_c82 bl_82 br_82 wl_71 vdd gnd cell_6t
Xbit_r72_c82 bl_82 br_82 wl_72 vdd gnd cell_6t
Xbit_r73_c82 bl_82 br_82 wl_73 vdd gnd cell_6t
Xbit_r74_c82 bl_82 br_82 wl_74 vdd gnd cell_6t
Xbit_r75_c82 bl_82 br_82 wl_75 vdd gnd cell_6t
Xbit_r76_c82 bl_82 br_82 wl_76 vdd gnd cell_6t
Xbit_r77_c82 bl_82 br_82 wl_77 vdd gnd cell_6t
Xbit_r78_c82 bl_82 br_82 wl_78 vdd gnd cell_6t
Xbit_r79_c82 bl_82 br_82 wl_79 vdd gnd cell_6t
Xbit_r80_c82 bl_82 br_82 wl_80 vdd gnd cell_6t
Xbit_r81_c82 bl_82 br_82 wl_81 vdd gnd cell_6t
Xbit_r82_c82 bl_82 br_82 wl_82 vdd gnd cell_6t
Xbit_r83_c82 bl_82 br_82 wl_83 vdd gnd cell_6t
Xbit_r84_c82 bl_82 br_82 wl_84 vdd gnd cell_6t
Xbit_r85_c82 bl_82 br_82 wl_85 vdd gnd cell_6t
Xbit_r86_c82 bl_82 br_82 wl_86 vdd gnd cell_6t
Xbit_r87_c82 bl_82 br_82 wl_87 vdd gnd cell_6t
Xbit_r88_c82 bl_82 br_82 wl_88 vdd gnd cell_6t
Xbit_r89_c82 bl_82 br_82 wl_89 vdd gnd cell_6t
Xbit_r90_c82 bl_82 br_82 wl_90 vdd gnd cell_6t
Xbit_r91_c82 bl_82 br_82 wl_91 vdd gnd cell_6t
Xbit_r92_c82 bl_82 br_82 wl_92 vdd gnd cell_6t
Xbit_r93_c82 bl_82 br_82 wl_93 vdd gnd cell_6t
Xbit_r94_c82 bl_82 br_82 wl_94 vdd gnd cell_6t
Xbit_r95_c82 bl_82 br_82 wl_95 vdd gnd cell_6t
Xbit_r96_c82 bl_82 br_82 wl_96 vdd gnd cell_6t
Xbit_r97_c82 bl_82 br_82 wl_97 vdd gnd cell_6t
Xbit_r98_c82 bl_82 br_82 wl_98 vdd gnd cell_6t
Xbit_r99_c82 bl_82 br_82 wl_99 vdd gnd cell_6t
Xbit_r100_c82 bl_82 br_82 wl_100 vdd gnd cell_6t
Xbit_r101_c82 bl_82 br_82 wl_101 vdd gnd cell_6t
Xbit_r102_c82 bl_82 br_82 wl_102 vdd gnd cell_6t
Xbit_r103_c82 bl_82 br_82 wl_103 vdd gnd cell_6t
Xbit_r104_c82 bl_82 br_82 wl_104 vdd gnd cell_6t
Xbit_r105_c82 bl_82 br_82 wl_105 vdd gnd cell_6t
Xbit_r106_c82 bl_82 br_82 wl_106 vdd gnd cell_6t
Xbit_r107_c82 bl_82 br_82 wl_107 vdd gnd cell_6t
Xbit_r108_c82 bl_82 br_82 wl_108 vdd gnd cell_6t
Xbit_r109_c82 bl_82 br_82 wl_109 vdd gnd cell_6t
Xbit_r110_c82 bl_82 br_82 wl_110 vdd gnd cell_6t
Xbit_r111_c82 bl_82 br_82 wl_111 vdd gnd cell_6t
Xbit_r112_c82 bl_82 br_82 wl_112 vdd gnd cell_6t
Xbit_r113_c82 bl_82 br_82 wl_113 vdd gnd cell_6t
Xbit_r114_c82 bl_82 br_82 wl_114 vdd gnd cell_6t
Xbit_r115_c82 bl_82 br_82 wl_115 vdd gnd cell_6t
Xbit_r116_c82 bl_82 br_82 wl_116 vdd gnd cell_6t
Xbit_r117_c82 bl_82 br_82 wl_117 vdd gnd cell_6t
Xbit_r118_c82 bl_82 br_82 wl_118 vdd gnd cell_6t
Xbit_r119_c82 bl_82 br_82 wl_119 vdd gnd cell_6t
Xbit_r120_c82 bl_82 br_82 wl_120 vdd gnd cell_6t
Xbit_r121_c82 bl_82 br_82 wl_121 vdd gnd cell_6t
Xbit_r122_c82 bl_82 br_82 wl_122 vdd gnd cell_6t
Xbit_r123_c82 bl_82 br_82 wl_123 vdd gnd cell_6t
Xbit_r124_c82 bl_82 br_82 wl_124 vdd gnd cell_6t
Xbit_r125_c82 bl_82 br_82 wl_125 vdd gnd cell_6t
Xbit_r126_c82 bl_82 br_82 wl_126 vdd gnd cell_6t
Xbit_r127_c82 bl_82 br_82 wl_127 vdd gnd cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd cell_6t
Xbit_r1_c83 bl_83 br_83 wl_1 vdd gnd cell_6t
Xbit_r2_c83 bl_83 br_83 wl_2 vdd gnd cell_6t
Xbit_r3_c83 bl_83 br_83 wl_3 vdd gnd cell_6t
Xbit_r4_c83 bl_83 br_83 wl_4 vdd gnd cell_6t
Xbit_r5_c83 bl_83 br_83 wl_5 vdd gnd cell_6t
Xbit_r6_c83 bl_83 br_83 wl_6 vdd gnd cell_6t
Xbit_r7_c83 bl_83 br_83 wl_7 vdd gnd cell_6t
Xbit_r8_c83 bl_83 br_83 wl_8 vdd gnd cell_6t
Xbit_r9_c83 bl_83 br_83 wl_9 vdd gnd cell_6t
Xbit_r10_c83 bl_83 br_83 wl_10 vdd gnd cell_6t
Xbit_r11_c83 bl_83 br_83 wl_11 vdd gnd cell_6t
Xbit_r12_c83 bl_83 br_83 wl_12 vdd gnd cell_6t
Xbit_r13_c83 bl_83 br_83 wl_13 vdd gnd cell_6t
Xbit_r14_c83 bl_83 br_83 wl_14 vdd gnd cell_6t
Xbit_r15_c83 bl_83 br_83 wl_15 vdd gnd cell_6t
Xbit_r16_c83 bl_83 br_83 wl_16 vdd gnd cell_6t
Xbit_r17_c83 bl_83 br_83 wl_17 vdd gnd cell_6t
Xbit_r18_c83 bl_83 br_83 wl_18 vdd gnd cell_6t
Xbit_r19_c83 bl_83 br_83 wl_19 vdd gnd cell_6t
Xbit_r20_c83 bl_83 br_83 wl_20 vdd gnd cell_6t
Xbit_r21_c83 bl_83 br_83 wl_21 vdd gnd cell_6t
Xbit_r22_c83 bl_83 br_83 wl_22 vdd gnd cell_6t
Xbit_r23_c83 bl_83 br_83 wl_23 vdd gnd cell_6t
Xbit_r24_c83 bl_83 br_83 wl_24 vdd gnd cell_6t
Xbit_r25_c83 bl_83 br_83 wl_25 vdd gnd cell_6t
Xbit_r26_c83 bl_83 br_83 wl_26 vdd gnd cell_6t
Xbit_r27_c83 bl_83 br_83 wl_27 vdd gnd cell_6t
Xbit_r28_c83 bl_83 br_83 wl_28 vdd gnd cell_6t
Xbit_r29_c83 bl_83 br_83 wl_29 vdd gnd cell_6t
Xbit_r30_c83 bl_83 br_83 wl_30 vdd gnd cell_6t
Xbit_r31_c83 bl_83 br_83 wl_31 vdd gnd cell_6t
Xbit_r32_c83 bl_83 br_83 wl_32 vdd gnd cell_6t
Xbit_r33_c83 bl_83 br_83 wl_33 vdd gnd cell_6t
Xbit_r34_c83 bl_83 br_83 wl_34 vdd gnd cell_6t
Xbit_r35_c83 bl_83 br_83 wl_35 vdd gnd cell_6t
Xbit_r36_c83 bl_83 br_83 wl_36 vdd gnd cell_6t
Xbit_r37_c83 bl_83 br_83 wl_37 vdd gnd cell_6t
Xbit_r38_c83 bl_83 br_83 wl_38 vdd gnd cell_6t
Xbit_r39_c83 bl_83 br_83 wl_39 vdd gnd cell_6t
Xbit_r40_c83 bl_83 br_83 wl_40 vdd gnd cell_6t
Xbit_r41_c83 bl_83 br_83 wl_41 vdd gnd cell_6t
Xbit_r42_c83 bl_83 br_83 wl_42 vdd gnd cell_6t
Xbit_r43_c83 bl_83 br_83 wl_43 vdd gnd cell_6t
Xbit_r44_c83 bl_83 br_83 wl_44 vdd gnd cell_6t
Xbit_r45_c83 bl_83 br_83 wl_45 vdd gnd cell_6t
Xbit_r46_c83 bl_83 br_83 wl_46 vdd gnd cell_6t
Xbit_r47_c83 bl_83 br_83 wl_47 vdd gnd cell_6t
Xbit_r48_c83 bl_83 br_83 wl_48 vdd gnd cell_6t
Xbit_r49_c83 bl_83 br_83 wl_49 vdd gnd cell_6t
Xbit_r50_c83 bl_83 br_83 wl_50 vdd gnd cell_6t
Xbit_r51_c83 bl_83 br_83 wl_51 vdd gnd cell_6t
Xbit_r52_c83 bl_83 br_83 wl_52 vdd gnd cell_6t
Xbit_r53_c83 bl_83 br_83 wl_53 vdd gnd cell_6t
Xbit_r54_c83 bl_83 br_83 wl_54 vdd gnd cell_6t
Xbit_r55_c83 bl_83 br_83 wl_55 vdd gnd cell_6t
Xbit_r56_c83 bl_83 br_83 wl_56 vdd gnd cell_6t
Xbit_r57_c83 bl_83 br_83 wl_57 vdd gnd cell_6t
Xbit_r58_c83 bl_83 br_83 wl_58 vdd gnd cell_6t
Xbit_r59_c83 bl_83 br_83 wl_59 vdd gnd cell_6t
Xbit_r60_c83 bl_83 br_83 wl_60 vdd gnd cell_6t
Xbit_r61_c83 bl_83 br_83 wl_61 vdd gnd cell_6t
Xbit_r62_c83 bl_83 br_83 wl_62 vdd gnd cell_6t
Xbit_r63_c83 bl_83 br_83 wl_63 vdd gnd cell_6t
Xbit_r64_c83 bl_83 br_83 wl_64 vdd gnd cell_6t
Xbit_r65_c83 bl_83 br_83 wl_65 vdd gnd cell_6t
Xbit_r66_c83 bl_83 br_83 wl_66 vdd gnd cell_6t
Xbit_r67_c83 bl_83 br_83 wl_67 vdd gnd cell_6t
Xbit_r68_c83 bl_83 br_83 wl_68 vdd gnd cell_6t
Xbit_r69_c83 bl_83 br_83 wl_69 vdd gnd cell_6t
Xbit_r70_c83 bl_83 br_83 wl_70 vdd gnd cell_6t
Xbit_r71_c83 bl_83 br_83 wl_71 vdd gnd cell_6t
Xbit_r72_c83 bl_83 br_83 wl_72 vdd gnd cell_6t
Xbit_r73_c83 bl_83 br_83 wl_73 vdd gnd cell_6t
Xbit_r74_c83 bl_83 br_83 wl_74 vdd gnd cell_6t
Xbit_r75_c83 bl_83 br_83 wl_75 vdd gnd cell_6t
Xbit_r76_c83 bl_83 br_83 wl_76 vdd gnd cell_6t
Xbit_r77_c83 bl_83 br_83 wl_77 vdd gnd cell_6t
Xbit_r78_c83 bl_83 br_83 wl_78 vdd gnd cell_6t
Xbit_r79_c83 bl_83 br_83 wl_79 vdd gnd cell_6t
Xbit_r80_c83 bl_83 br_83 wl_80 vdd gnd cell_6t
Xbit_r81_c83 bl_83 br_83 wl_81 vdd gnd cell_6t
Xbit_r82_c83 bl_83 br_83 wl_82 vdd gnd cell_6t
Xbit_r83_c83 bl_83 br_83 wl_83 vdd gnd cell_6t
Xbit_r84_c83 bl_83 br_83 wl_84 vdd gnd cell_6t
Xbit_r85_c83 bl_83 br_83 wl_85 vdd gnd cell_6t
Xbit_r86_c83 bl_83 br_83 wl_86 vdd gnd cell_6t
Xbit_r87_c83 bl_83 br_83 wl_87 vdd gnd cell_6t
Xbit_r88_c83 bl_83 br_83 wl_88 vdd gnd cell_6t
Xbit_r89_c83 bl_83 br_83 wl_89 vdd gnd cell_6t
Xbit_r90_c83 bl_83 br_83 wl_90 vdd gnd cell_6t
Xbit_r91_c83 bl_83 br_83 wl_91 vdd gnd cell_6t
Xbit_r92_c83 bl_83 br_83 wl_92 vdd gnd cell_6t
Xbit_r93_c83 bl_83 br_83 wl_93 vdd gnd cell_6t
Xbit_r94_c83 bl_83 br_83 wl_94 vdd gnd cell_6t
Xbit_r95_c83 bl_83 br_83 wl_95 vdd gnd cell_6t
Xbit_r96_c83 bl_83 br_83 wl_96 vdd gnd cell_6t
Xbit_r97_c83 bl_83 br_83 wl_97 vdd gnd cell_6t
Xbit_r98_c83 bl_83 br_83 wl_98 vdd gnd cell_6t
Xbit_r99_c83 bl_83 br_83 wl_99 vdd gnd cell_6t
Xbit_r100_c83 bl_83 br_83 wl_100 vdd gnd cell_6t
Xbit_r101_c83 bl_83 br_83 wl_101 vdd gnd cell_6t
Xbit_r102_c83 bl_83 br_83 wl_102 vdd gnd cell_6t
Xbit_r103_c83 bl_83 br_83 wl_103 vdd gnd cell_6t
Xbit_r104_c83 bl_83 br_83 wl_104 vdd gnd cell_6t
Xbit_r105_c83 bl_83 br_83 wl_105 vdd gnd cell_6t
Xbit_r106_c83 bl_83 br_83 wl_106 vdd gnd cell_6t
Xbit_r107_c83 bl_83 br_83 wl_107 vdd gnd cell_6t
Xbit_r108_c83 bl_83 br_83 wl_108 vdd gnd cell_6t
Xbit_r109_c83 bl_83 br_83 wl_109 vdd gnd cell_6t
Xbit_r110_c83 bl_83 br_83 wl_110 vdd gnd cell_6t
Xbit_r111_c83 bl_83 br_83 wl_111 vdd gnd cell_6t
Xbit_r112_c83 bl_83 br_83 wl_112 vdd gnd cell_6t
Xbit_r113_c83 bl_83 br_83 wl_113 vdd gnd cell_6t
Xbit_r114_c83 bl_83 br_83 wl_114 vdd gnd cell_6t
Xbit_r115_c83 bl_83 br_83 wl_115 vdd gnd cell_6t
Xbit_r116_c83 bl_83 br_83 wl_116 vdd gnd cell_6t
Xbit_r117_c83 bl_83 br_83 wl_117 vdd gnd cell_6t
Xbit_r118_c83 bl_83 br_83 wl_118 vdd gnd cell_6t
Xbit_r119_c83 bl_83 br_83 wl_119 vdd gnd cell_6t
Xbit_r120_c83 bl_83 br_83 wl_120 vdd gnd cell_6t
Xbit_r121_c83 bl_83 br_83 wl_121 vdd gnd cell_6t
Xbit_r122_c83 bl_83 br_83 wl_122 vdd gnd cell_6t
Xbit_r123_c83 bl_83 br_83 wl_123 vdd gnd cell_6t
Xbit_r124_c83 bl_83 br_83 wl_124 vdd gnd cell_6t
Xbit_r125_c83 bl_83 br_83 wl_125 vdd gnd cell_6t
Xbit_r126_c83 bl_83 br_83 wl_126 vdd gnd cell_6t
Xbit_r127_c83 bl_83 br_83 wl_127 vdd gnd cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd cell_6t
Xbit_r1_c84 bl_84 br_84 wl_1 vdd gnd cell_6t
Xbit_r2_c84 bl_84 br_84 wl_2 vdd gnd cell_6t
Xbit_r3_c84 bl_84 br_84 wl_3 vdd gnd cell_6t
Xbit_r4_c84 bl_84 br_84 wl_4 vdd gnd cell_6t
Xbit_r5_c84 bl_84 br_84 wl_5 vdd gnd cell_6t
Xbit_r6_c84 bl_84 br_84 wl_6 vdd gnd cell_6t
Xbit_r7_c84 bl_84 br_84 wl_7 vdd gnd cell_6t
Xbit_r8_c84 bl_84 br_84 wl_8 vdd gnd cell_6t
Xbit_r9_c84 bl_84 br_84 wl_9 vdd gnd cell_6t
Xbit_r10_c84 bl_84 br_84 wl_10 vdd gnd cell_6t
Xbit_r11_c84 bl_84 br_84 wl_11 vdd gnd cell_6t
Xbit_r12_c84 bl_84 br_84 wl_12 vdd gnd cell_6t
Xbit_r13_c84 bl_84 br_84 wl_13 vdd gnd cell_6t
Xbit_r14_c84 bl_84 br_84 wl_14 vdd gnd cell_6t
Xbit_r15_c84 bl_84 br_84 wl_15 vdd gnd cell_6t
Xbit_r16_c84 bl_84 br_84 wl_16 vdd gnd cell_6t
Xbit_r17_c84 bl_84 br_84 wl_17 vdd gnd cell_6t
Xbit_r18_c84 bl_84 br_84 wl_18 vdd gnd cell_6t
Xbit_r19_c84 bl_84 br_84 wl_19 vdd gnd cell_6t
Xbit_r20_c84 bl_84 br_84 wl_20 vdd gnd cell_6t
Xbit_r21_c84 bl_84 br_84 wl_21 vdd gnd cell_6t
Xbit_r22_c84 bl_84 br_84 wl_22 vdd gnd cell_6t
Xbit_r23_c84 bl_84 br_84 wl_23 vdd gnd cell_6t
Xbit_r24_c84 bl_84 br_84 wl_24 vdd gnd cell_6t
Xbit_r25_c84 bl_84 br_84 wl_25 vdd gnd cell_6t
Xbit_r26_c84 bl_84 br_84 wl_26 vdd gnd cell_6t
Xbit_r27_c84 bl_84 br_84 wl_27 vdd gnd cell_6t
Xbit_r28_c84 bl_84 br_84 wl_28 vdd gnd cell_6t
Xbit_r29_c84 bl_84 br_84 wl_29 vdd gnd cell_6t
Xbit_r30_c84 bl_84 br_84 wl_30 vdd gnd cell_6t
Xbit_r31_c84 bl_84 br_84 wl_31 vdd gnd cell_6t
Xbit_r32_c84 bl_84 br_84 wl_32 vdd gnd cell_6t
Xbit_r33_c84 bl_84 br_84 wl_33 vdd gnd cell_6t
Xbit_r34_c84 bl_84 br_84 wl_34 vdd gnd cell_6t
Xbit_r35_c84 bl_84 br_84 wl_35 vdd gnd cell_6t
Xbit_r36_c84 bl_84 br_84 wl_36 vdd gnd cell_6t
Xbit_r37_c84 bl_84 br_84 wl_37 vdd gnd cell_6t
Xbit_r38_c84 bl_84 br_84 wl_38 vdd gnd cell_6t
Xbit_r39_c84 bl_84 br_84 wl_39 vdd gnd cell_6t
Xbit_r40_c84 bl_84 br_84 wl_40 vdd gnd cell_6t
Xbit_r41_c84 bl_84 br_84 wl_41 vdd gnd cell_6t
Xbit_r42_c84 bl_84 br_84 wl_42 vdd gnd cell_6t
Xbit_r43_c84 bl_84 br_84 wl_43 vdd gnd cell_6t
Xbit_r44_c84 bl_84 br_84 wl_44 vdd gnd cell_6t
Xbit_r45_c84 bl_84 br_84 wl_45 vdd gnd cell_6t
Xbit_r46_c84 bl_84 br_84 wl_46 vdd gnd cell_6t
Xbit_r47_c84 bl_84 br_84 wl_47 vdd gnd cell_6t
Xbit_r48_c84 bl_84 br_84 wl_48 vdd gnd cell_6t
Xbit_r49_c84 bl_84 br_84 wl_49 vdd gnd cell_6t
Xbit_r50_c84 bl_84 br_84 wl_50 vdd gnd cell_6t
Xbit_r51_c84 bl_84 br_84 wl_51 vdd gnd cell_6t
Xbit_r52_c84 bl_84 br_84 wl_52 vdd gnd cell_6t
Xbit_r53_c84 bl_84 br_84 wl_53 vdd gnd cell_6t
Xbit_r54_c84 bl_84 br_84 wl_54 vdd gnd cell_6t
Xbit_r55_c84 bl_84 br_84 wl_55 vdd gnd cell_6t
Xbit_r56_c84 bl_84 br_84 wl_56 vdd gnd cell_6t
Xbit_r57_c84 bl_84 br_84 wl_57 vdd gnd cell_6t
Xbit_r58_c84 bl_84 br_84 wl_58 vdd gnd cell_6t
Xbit_r59_c84 bl_84 br_84 wl_59 vdd gnd cell_6t
Xbit_r60_c84 bl_84 br_84 wl_60 vdd gnd cell_6t
Xbit_r61_c84 bl_84 br_84 wl_61 vdd gnd cell_6t
Xbit_r62_c84 bl_84 br_84 wl_62 vdd gnd cell_6t
Xbit_r63_c84 bl_84 br_84 wl_63 vdd gnd cell_6t
Xbit_r64_c84 bl_84 br_84 wl_64 vdd gnd cell_6t
Xbit_r65_c84 bl_84 br_84 wl_65 vdd gnd cell_6t
Xbit_r66_c84 bl_84 br_84 wl_66 vdd gnd cell_6t
Xbit_r67_c84 bl_84 br_84 wl_67 vdd gnd cell_6t
Xbit_r68_c84 bl_84 br_84 wl_68 vdd gnd cell_6t
Xbit_r69_c84 bl_84 br_84 wl_69 vdd gnd cell_6t
Xbit_r70_c84 bl_84 br_84 wl_70 vdd gnd cell_6t
Xbit_r71_c84 bl_84 br_84 wl_71 vdd gnd cell_6t
Xbit_r72_c84 bl_84 br_84 wl_72 vdd gnd cell_6t
Xbit_r73_c84 bl_84 br_84 wl_73 vdd gnd cell_6t
Xbit_r74_c84 bl_84 br_84 wl_74 vdd gnd cell_6t
Xbit_r75_c84 bl_84 br_84 wl_75 vdd gnd cell_6t
Xbit_r76_c84 bl_84 br_84 wl_76 vdd gnd cell_6t
Xbit_r77_c84 bl_84 br_84 wl_77 vdd gnd cell_6t
Xbit_r78_c84 bl_84 br_84 wl_78 vdd gnd cell_6t
Xbit_r79_c84 bl_84 br_84 wl_79 vdd gnd cell_6t
Xbit_r80_c84 bl_84 br_84 wl_80 vdd gnd cell_6t
Xbit_r81_c84 bl_84 br_84 wl_81 vdd gnd cell_6t
Xbit_r82_c84 bl_84 br_84 wl_82 vdd gnd cell_6t
Xbit_r83_c84 bl_84 br_84 wl_83 vdd gnd cell_6t
Xbit_r84_c84 bl_84 br_84 wl_84 vdd gnd cell_6t
Xbit_r85_c84 bl_84 br_84 wl_85 vdd gnd cell_6t
Xbit_r86_c84 bl_84 br_84 wl_86 vdd gnd cell_6t
Xbit_r87_c84 bl_84 br_84 wl_87 vdd gnd cell_6t
Xbit_r88_c84 bl_84 br_84 wl_88 vdd gnd cell_6t
Xbit_r89_c84 bl_84 br_84 wl_89 vdd gnd cell_6t
Xbit_r90_c84 bl_84 br_84 wl_90 vdd gnd cell_6t
Xbit_r91_c84 bl_84 br_84 wl_91 vdd gnd cell_6t
Xbit_r92_c84 bl_84 br_84 wl_92 vdd gnd cell_6t
Xbit_r93_c84 bl_84 br_84 wl_93 vdd gnd cell_6t
Xbit_r94_c84 bl_84 br_84 wl_94 vdd gnd cell_6t
Xbit_r95_c84 bl_84 br_84 wl_95 vdd gnd cell_6t
Xbit_r96_c84 bl_84 br_84 wl_96 vdd gnd cell_6t
Xbit_r97_c84 bl_84 br_84 wl_97 vdd gnd cell_6t
Xbit_r98_c84 bl_84 br_84 wl_98 vdd gnd cell_6t
Xbit_r99_c84 bl_84 br_84 wl_99 vdd gnd cell_6t
Xbit_r100_c84 bl_84 br_84 wl_100 vdd gnd cell_6t
Xbit_r101_c84 bl_84 br_84 wl_101 vdd gnd cell_6t
Xbit_r102_c84 bl_84 br_84 wl_102 vdd gnd cell_6t
Xbit_r103_c84 bl_84 br_84 wl_103 vdd gnd cell_6t
Xbit_r104_c84 bl_84 br_84 wl_104 vdd gnd cell_6t
Xbit_r105_c84 bl_84 br_84 wl_105 vdd gnd cell_6t
Xbit_r106_c84 bl_84 br_84 wl_106 vdd gnd cell_6t
Xbit_r107_c84 bl_84 br_84 wl_107 vdd gnd cell_6t
Xbit_r108_c84 bl_84 br_84 wl_108 vdd gnd cell_6t
Xbit_r109_c84 bl_84 br_84 wl_109 vdd gnd cell_6t
Xbit_r110_c84 bl_84 br_84 wl_110 vdd gnd cell_6t
Xbit_r111_c84 bl_84 br_84 wl_111 vdd gnd cell_6t
Xbit_r112_c84 bl_84 br_84 wl_112 vdd gnd cell_6t
Xbit_r113_c84 bl_84 br_84 wl_113 vdd gnd cell_6t
Xbit_r114_c84 bl_84 br_84 wl_114 vdd gnd cell_6t
Xbit_r115_c84 bl_84 br_84 wl_115 vdd gnd cell_6t
Xbit_r116_c84 bl_84 br_84 wl_116 vdd gnd cell_6t
Xbit_r117_c84 bl_84 br_84 wl_117 vdd gnd cell_6t
Xbit_r118_c84 bl_84 br_84 wl_118 vdd gnd cell_6t
Xbit_r119_c84 bl_84 br_84 wl_119 vdd gnd cell_6t
Xbit_r120_c84 bl_84 br_84 wl_120 vdd gnd cell_6t
Xbit_r121_c84 bl_84 br_84 wl_121 vdd gnd cell_6t
Xbit_r122_c84 bl_84 br_84 wl_122 vdd gnd cell_6t
Xbit_r123_c84 bl_84 br_84 wl_123 vdd gnd cell_6t
Xbit_r124_c84 bl_84 br_84 wl_124 vdd gnd cell_6t
Xbit_r125_c84 bl_84 br_84 wl_125 vdd gnd cell_6t
Xbit_r126_c84 bl_84 br_84 wl_126 vdd gnd cell_6t
Xbit_r127_c84 bl_84 br_84 wl_127 vdd gnd cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd cell_6t
Xbit_r1_c85 bl_85 br_85 wl_1 vdd gnd cell_6t
Xbit_r2_c85 bl_85 br_85 wl_2 vdd gnd cell_6t
Xbit_r3_c85 bl_85 br_85 wl_3 vdd gnd cell_6t
Xbit_r4_c85 bl_85 br_85 wl_4 vdd gnd cell_6t
Xbit_r5_c85 bl_85 br_85 wl_5 vdd gnd cell_6t
Xbit_r6_c85 bl_85 br_85 wl_6 vdd gnd cell_6t
Xbit_r7_c85 bl_85 br_85 wl_7 vdd gnd cell_6t
Xbit_r8_c85 bl_85 br_85 wl_8 vdd gnd cell_6t
Xbit_r9_c85 bl_85 br_85 wl_9 vdd gnd cell_6t
Xbit_r10_c85 bl_85 br_85 wl_10 vdd gnd cell_6t
Xbit_r11_c85 bl_85 br_85 wl_11 vdd gnd cell_6t
Xbit_r12_c85 bl_85 br_85 wl_12 vdd gnd cell_6t
Xbit_r13_c85 bl_85 br_85 wl_13 vdd gnd cell_6t
Xbit_r14_c85 bl_85 br_85 wl_14 vdd gnd cell_6t
Xbit_r15_c85 bl_85 br_85 wl_15 vdd gnd cell_6t
Xbit_r16_c85 bl_85 br_85 wl_16 vdd gnd cell_6t
Xbit_r17_c85 bl_85 br_85 wl_17 vdd gnd cell_6t
Xbit_r18_c85 bl_85 br_85 wl_18 vdd gnd cell_6t
Xbit_r19_c85 bl_85 br_85 wl_19 vdd gnd cell_6t
Xbit_r20_c85 bl_85 br_85 wl_20 vdd gnd cell_6t
Xbit_r21_c85 bl_85 br_85 wl_21 vdd gnd cell_6t
Xbit_r22_c85 bl_85 br_85 wl_22 vdd gnd cell_6t
Xbit_r23_c85 bl_85 br_85 wl_23 vdd gnd cell_6t
Xbit_r24_c85 bl_85 br_85 wl_24 vdd gnd cell_6t
Xbit_r25_c85 bl_85 br_85 wl_25 vdd gnd cell_6t
Xbit_r26_c85 bl_85 br_85 wl_26 vdd gnd cell_6t
Xbit_r27_c85 bl_85 br_85 wl_27 vdd gnd cell_6t
Xbit_r28_c85 bl_85 br_85 wl_28 vdd gnd cell_6t
Xbit_r29_c85 bl_85 br_85 wl_29 vdd gnd cell_6t
Xbit_r30_c85 bl_85 br_85 wl_30 vdd gnd cell_6t
Xbit_r31_c85 bl_85 br_85 wl_31 vdd gnd cell_6t
Xbit_r32_c85 bl_85 br_85 wl_32 vdd gnd cell_6t
Xbit_r33_c85 bl_85 br_85 wl_33 vdd gnd cell_6t
Xbit_r34_c85 bl_85 br_85 wl_34 vdd gnd cell_6t
Xbit_r35_c85 bl_85 br_85 wl_35 vdd gnd cell_6t
Xbit_r36_c85 bl_85 br_85 wl_36 vdd gnd cell_6t
Xbit_r37_c85 bl_85 br_85 wl_37 vdd gnd cell_6t
Xbit_r38_c85 bl_85 br_85 wl_38 vdd gnd cell_6t
Xbit_r39_c85 bl_85 br_85 wl_39 vdd gnd cell_6t
Xbit_r40_c85 bl_85 br_85 wl_40 vdd gnd cell_6t
Xbit_r41_c85 bl_85 br_85 wl_41 vdd gnd cell_6t
Xbit_r42_c85 bl_85 br_85 wl_42 vdd gnd cell_6t
Xbit_r43_c85 bl_85 br_85 wl_43 vdd gnd cell_6t
Xbit_r44_c85 bl_85 br_85 wl_44 vdd gnd cell_6t
Xbit_r45_c85 bl_85 br_85 wl_45 vdd gnd cell_6t
Xbit_r46_c85 bl_85 br_85 wl_46 vdd gnd cell_6t
Xbit_r47_c85 bl_85 br_85 wl_47 vdd gnd cell_6t
Xbit_r48_c85 bl_85 br_85 wl_48 vdd gnd cell_6t
Xbit_r49_c85 bl_85 br_85 wl_49 vdd gnd cell_6t
Xbit_r50_c85 bl_85 br_85 wl_50 vdd gnd cell_6t
Xbit_r51_c85 bl_85 br_85 wl_51 vdd gnd cell_6t
Xbit_r52_c85 bl_85 br_85 wl_52 vdd gnd cell_6t
Xbit_r53_c85 bl_85 br_85 wl_53 vdd gnd cell_6t
Xbit_r54_c85 bl_85 br_85 wl_54 vdd gnd cell_6t
Xbit_r55_c85 bl_85 br_85 wl_55 vdd gnd cell_6t
Xbit_r56_c85 bl_85 br_85 wl_56 vdd gnd cell_6t
Xbit_r57_c85 bl_85 br_85 wl_57 vdd gnd cell_6t
Xbit_r58_c85 bl_85 br_85 wl_58 vdd gnd cell_6t
Xbit_r59_c85 bl_85 br_85 wl_59 vdd gnd cell_6t
Xbit_r60_c85 bl_85 br_85 wl_60 vdd gnd cell_6t
Xbit_r61_c85 bl_85 br_85 wl_61 vdd gnd cell_6t
Xbit_r62_c85 bl_85 br_85 wl_62 vdd gnd cell_6t
Xbit_r63_c85 bl_85 br_85 wl_63 vdd gnd cell_6t
Xbit_r64_c85 bl_85 br_85 wl_64 vdd gnd cell_6t
Xbit_r65_c85 bl_85 br_85 wl_65 vdd gnd cell_6t
Xbit_r66_c85 bl_85 br_85 wl_66 vdd gnd cell_6t
Xbit_r67_c85 bl_85 br_85 wl_67 vdd gnd cell_6t
Xbit_r68_c85 bl_85 br_85 wl_68 vdd gnd cell_6t
Xbit_r69_c85 bl_85 br_85 wl_69 vdd gnd cell_6t
Xbit_r70_c85 bl_85 br_85 wl_70 vdd gnd cell_6t
Xbit_r71_c85 bl_85 br_85 wl_71 vdd gnd cell_6t
Xbit_r72_c85 bl_85 br_85 wl_72 vdd gnd cell_6t
Xbit_r73_c85 bl_85 br_85 wl_73 vdd gnd cell_6t
Xbit_r74_c85 bl_85 br_85 wl_74 vdd gnd cell_6t
Xbit_r75_c85 bl_85 br_85 wl_75 vdd gnd cell_6t
Xbit_r76_c85 bl_85 br_85 wl_76 vdd gnd cell_6t
Xbit_r77_c85 bl_85 br_85 wl_77 vdd gnd cell_6t
Xbit_r78_c85 bl_85 br_85 wl_78 vdd gnd cell_6t
Xbit_r79_c85 bl_85 br_85 wl_79 vdd gnd cell_6t
Xbit_r80_c85 bl_85 br_85 wl_80 vdd gnd cell_6t
Xbit_r81_c85 bl_85 br_85 wl_81 vdd gnd cell_6t
Xbit_r82_c85 bl_85 br_85 wl_82 vdd gnd cell_6t
Xbit_r83_c85 bl_85 br_85 wl_83 vdd gnd cell_6t
Xbit_r84_c85 bl_85 br_85 wl_84 vdd gnd cell_6t
Xbit_r85_c85 bl_85 br_85 wl_85 vdd gnd cell_6t
Xbit_r86_c85 bl_85 br_85 wl_86 vdd gnd cell_6t
Xbit_r87_c85 bl_85 br_85 wl_87 vdd gnd cell_6t
Xbit_r88_c85 bl_85 br_85 wl_88 vdd gnd cell_6t
Xbit_r89_c85 bl_85 br_85 wl_89 vdd gnd cell_6t
Xbit_r90_c85 bl_85 br_85 wl_90 vdd gnd cell_6t
Xbit_r91_c85 bl_85 br_85 wl_91 vdd gnd cell_6t
Xbit_r92_c85 bl_85 br_85 wl_92 vdd gnd cell_6t
Xbit_r93_c85 bl_85 br_85 wl_93 vdd gnd cell_6t
Xbit_r94_c85 bl_85 br_85 wl_94 vdd gnd cell_6t
Xbit_r95_c85 bl_85 br_85 wl_95 vdd gnd cell_6t
Xbit_r96_c85 bl_85 br_85 wl_96 vdd gnd cell_6t
Xbit_r97_c85 bl_85 br_85 wl_97 vdd gnd cell_6t
Xbit_r98_c85 bl_85 br_85 wl_98 vdd gnd cell_6t
Xbit_r99_c85 bl_85 br_85 wl_99 vdd gnd cell_6t
Xbit_r100_c85 bl_85 br_85 wl_100 vdd gnd cell_6t
Xbit_r101_c85 bl_85 br_85 wl_101 vdd gnd cell_6t
Xbit_r102_c85 bl_85 br_85 wl_102 vdd gnd cell_6t
Xbit_r103_c85 bl_85 br_85 wl_103 vdd gnd cell_6t
Xbit_r104_c85 bl_85 br_85 wl_104 vdd gnd cell_6t
Xbit_r105_c85 bl_85 br_85 wl_105 vdd gnd cell_6t
Xbit_r106_c85 bl_85 br_85 wl_106 vdd gnd cell_6t
Xbit_r107_c85 bl_85 br_85 wl_107 vdd gnd cell_6t
Xbit_r108_c85 bl_85 br_85 wl_108 vdd gnd cell_6t
Xbit_r109_c85 bl_85 br_85 wl_109 vdd gnd cell_6t
Xbit_r110_c85 bl_85 br_85 wl_110 vdd gnd cell_6t
Xbit_r111_c85 bl_85 br_85 wl_111 vdd gnd cell_6t
Xbit_r112_c85 bl_85 br_85 wl_112 vdd gnd cell_6t
Xbit_r113_c85 bl_85 br_85 wl_113 vdd gnd cell_6t
Xbit_r114_c85 bl_85 br_85 wl_114 vdd gnd cell_6t
Xbit_r115_c85 bl_85 br_85 wl_115 vdd gnd cell_6t
Xbit_r116_c85 bl_85 br_85 wl_116 vdd gnd cell_6t
Xbit_r117_c85 bl_85 br_85 wl_117 vdd gnd cell_6t
Xbit_r118_c85 bl_85 br_85 wl_118 vdd gnd cell_6t
Xbit_r119_c85 bl_85 br_85 wl_119 vdd gnd cell_6t
Xbit_r120_c85 bl_85 br_85 wl_120 vdd gnd cell_6t
Xbit_r121_c85 bl_85 br_85 wl_121 vdd gnd cell_6t
Xbit_r122_c85 bl_85 br_85 wl_122 vdd gnd cell_6t
Xbit_r123_c85 bl_85 br_85 wl_123 vdd gnd cell_6t
Xbit_r124_c85 bl_85 br_85 wl_124 vdd gnd cell_6t
Xbit_r125_c85 bl_85 br_85 wl_125 vdd gnd cell_6t
Xbit_r126_c85 bl_85 br_85 wl_126 vdd gnd cell_6t
Xbit_r127_c85 bl_85 br_85 wl_127 vdd gnd cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd cell_6t
Xbit_r1_c86 bl_86 br_86 wl_1 vdd gnd cell_6t
Xbit_r2_c86 bl_86 br_86 wl_2 vdd gnd cell_6t
Xbit_r3_c86 bl_86 br_86 wl_3 vdd gnd cell_6t
Xbit_r4_c86 bl_86 br_86 wl_4 vdd gnd cell_6t
Xbit_r5_c86 bl_86 br_86 wl_5 vdd gnd cell_6t
Xbit_r6_c86 bl_86 br_86 wl_6 vdd gnd cell_6t
Xbit_r7_c86 bl_86 br_86 wl_7 vdd gnd cell_6t
Xbit_r8_c86 bl_86 br_86 wl_8 vdd gnd cell_6t
Xbit_r9_c86 bl_86 br_86 wl_9 vdd gnd cell_6t
Xbit_r10_c86 bl_86 br_86 wl_10 vdd gnd cell_6t
Xbit_r11_c86 bl_86 br_86 wl_11 vdd gnd cell_6t
Xbit_r12_c86 bl_86 br_86 wl_12 vdd gnd cell_6t
Xbit_r13_c86 bl_86 br_86 wl_13 vdd gnd cell_6t
Xbit_r14_c86 bl_86 br_86 wl_14 vdd gnd cell_6t
Xbit_r15_c86 bl_86 br_86 wl_15 vdd gnd cell_6t
Xbit_r16_c86 bl_86 br_86 wl_16 vdd gnd cell_6t
Xbit_r17_c86 bl_86 br_86 wl_17 vdd gnd cell_6t
Xbit_r18_c86 bl_86 br_86 wl_18 vdd gnd cell_6t
Xbit_r19_c86 bl_86 br_86 wl_19 vdd gnd cell_6t
Xbit_r20_c86 bl_86 br_86 wl_20 vdd gnd cell_6t
Xbit_r21_c86 bl_86 br_86 wl_21 vdd gnd cell_6t
Xbit_r22_c86 bl_86 br_86 wl_22 vdd gnd cell_6t
Xbit_r23_c86 bl_86 br_86 wl_23 vdd gnd cell_6t
Xbit_r24_c86 bl_86 br_86 wl_24 vdd gnd cell_6t
Xbit_r25_c86 bl_86 br_86 wl_25 vdd gnd cell_6t
Xbit_r26_c86 bl_86 br_86 wl_26 vdd gnd cell_6t
Xbit_r27_c86 bl_86 br_86 wl_27 vdd gnd cell_6t
Xbit_r28_c86 bl_86 br_86 wl_28 vdd gnd cell_6t
Xbit_r29_c86 bl_86 br_86 wl_29 vdd gnd cell_6t
Xbit_r30_c86 bl_86 br_86 wl_30 vdd gnd cell_6t
Xbit_r31_c86 bl_86 br_86 wl_31 vdd gnd cell_6t
Xbit_r32_c86 bl_86 br_86 wl_32 vdd gnd cell_6t
Xbit_r33_c86 bl_86 br_86 wl_33 vdd gnd cell_6t
Xbit_r34_c86 bl_86 br_86 wl_34 vdd gnd cell_6t
Xbit_r35_c86 bl_86 br_86 wl_35 vdd gnd cell_6t
Xbit_r36_c86 bl_86 br_86 wl_36 vdd gnd cell_6t
Xbit_r37_c86 bl_86 br_86 wl_37 vdd gnd cell_6t
Xbit_r38_c86 bl_86 br_86 wl_38 vdd gnd cell_6t
Xbit_r39_c86 bl_86 br_86 wl_39 vdd gnd cell_6t
Xbit_r40_c86 bl_86 br_86 wl_40 vdd gnd cell_6t
Xbit_r41_c86 bl_86 br_86 wl_41 vdd gnd cell_6t
Xbit_r42_c86 bl_86 br_86 wl_42 vdd gnd cell_6t
Xbit_r43_c86 bl_86 br_86 wl_43 vdd gnd cell_6t
Xbit_r44_c86 bl_86 br_86 wl_44 vdd gnd cell_6t
Xbit_r45_c86 bl_86 br_86 wl_45 vdd gnd cell_6t
Xbit_r46_c86 bl_86 br_86 wl_46 vdd gnd cell_6t
Xbit_r47_c86 bl_86 br_86 wl_47 vdd gnd cell_6t
Xbit_r48_c86 bl_86 br_86 wl_48 vdd gnd cell_6t
Xbit_r49_c86 bl_86 br_86 wl_49 vdd gnd cell_6t
Xbit_r50_c86 bl_86 br_86 wl_50 vdd gnd cell_6t
Xbit_r51_c86 bl_86 br_86 wl_51 vdd gnd cell_6t
Xbit_r52_c86 bl_86 br_86 wl_52 vdd gnd cell_6t
Xbit_r53_c86 bl_86 br_86 wl_53 vdd gnd cell_6t
Xbit_r54_c86 bl_86 br_86 wl_54 vdd gnd cell_6t
Xbit_r55_c86 bl_86 br_86 wl_55 vdd gnd cell_6t
Xbit_r56_c86 bl_86 br_86 wl_56 vdd gnd cell_6t
Xbit_r57_c86 bl_86 br_86 wl_57 vdd gnd cell_6t
Xbit_r58_c86 bl_86 br_86 wl_58 vdd gnd cell_6t
Xbit_r59_c86 bl_86 br_86 wl_59 vdd gnd cell_6t
Xbit_r60_c86 bl_86 br_86 wl_60 vdd gnd cell_6t
Xbit_r61_c86 bl_86 br_86 wl_61 vdd gnd cell_6t
Xbit_r62_c86 bl_86 br_86 wl_62 vdd gnd cell_6t
Xbit_r63_c86 bl_86 br_86 wl_63 vdd gnd cell_6t
Xbit_r64_c86 bl_86 br_86 wl_64 vdd gnd cell_6t
Xbit_r65_c86 bl_86 br_86 wl_65 vdd gnd cell_6t
Xbit_r66_c86 bl_86 br_86 wl_66 vdd gnd cell_6t
Xbit_r67_c86 bl_86 br_86 wl_67 vdd gnd cell_6t
Xbit_r68_c86 bl_86 br_86 wl_68 vdd gnd cell_6t
Xbit_r69_c86 bl_86 br_86 wl_69 vdd gnd cell_6t
Xbit_r70_c86 bl_86 br_86 wl_70 vdd gnd cell_6t
Xbit_r71_c86 bl_86 br_86 wl_71 vdd gnd cell_6t
Xbit_r72_c86 bl_86 br_86 wl_72 vdd gnd cell_6t
Xbit_r73_c86 bl_86 br_86 wl_73 vdd gnd cell_6t
Xbit_r74_c86 bl_86 br_86 wl_74 vdd gnd cell_6t
Xbit_r75_c86 bl_86 br_86 wl_75 vdd gnd cell_6t
Xbit_r76_c86 bl_86 br_86 wl_76 vdd gnd cell_6t
Xbit_r77_c86 bl_86 br_86 wl_77 vdd gnd cell_6t
Xbit_r78_c86 bl_86 br_86 wl_78 vdd gnd cell_6t
Xbit_r79_c86 bl_86 br_86 wl_79 vdd gnd cell_6t
Xbit_r80_c86 bl_86 br_86 wl_80 vdd gnd cell_6t
Xbit_r81_c86 bl_86 br_86 wl_81 vdd gnd cell_6t
Xbit_r82_c86 bl_86 br_86 wl_82 vdd gnd cell_6t
Xbit_r83_c86 bl_86 br_86 wl_83 vdd gnd cell_6t
Xbit_r84_c86 bl_86 br_86 wl_84 vdd gnd cell_6t
Xbit_r85_c86 bl_86 br_86 wl_85 vdd gnd cell_6t
Xbit_r86_c86 bl_86 br_86 wl_86 vdd gnd cell_6t
Xbit_r87_c86 bl_86 br_86 wl_87 vdd gnd cell_6t
Xbit_r88_c86 bl_86 br_86 wl_88 vdd gnd cell_6t
Xbit_r89_c86 bl_86 br_86 wl_89 vdd gnd cell_6t
Xbit_r90_c86 bl_86 br_86 wl_90 vdd gnd cell_6t
Xbit_r91_c86 bl_86 br_86 wl_91 vdd gnd cell_6t
Xbit_r92_c86 bl_86 br_86 wl_92 vdd gnd cell_6t
Xbit_r93_c86 bl_86 br_86 wl_93 vdd gnd cell_6t
Xbit_r94_c86 bl_86 br_86 wl_94 vdd gnd cell_6t
Xbit_r95_c86 bl_86 br_86 wl_95 vdd gnd cell_6t
Xbit_r96_c86 bl_86 br_86 wl_96 vdd gnd cell_6t
Xbit_r97_c86 bl_86 br_86 wl_97 vdd gnd cell_6t
Xbit_r98_c86 bl_86 br_86 wl_98 vdd gnd cell_6t
Xbit_r99_c86 bl_86 br_86 wl_99 vdd gnd cell_6t
Xbit_r100_c86 bl_86 br_86 wl_100 vdd gnd cell_6t
Xbit_r101_c86 bl_86 br_86 wl_101 vdd gnd cell_6t
Xbit_r102_c86 bl_86 br_86 wl_102 vdd gnd cell_6t
Xbit_r103_c86 bl_86 br_86 wl_103 vdd gnd cell_6t
Xbit_r104_c86 bl_86 br_86 wl_104 vdd gnd cell_6t
Xbit_r105_c86 bl_86 br_86 wl_105 vdd gnd cell_6t
Xbit_r106_c86 bl_86 br_86 wl_106 vdd gnd cell_6t
Xbit_r107_c86 bl_86 br_86 wl_107 vdd gnd cell_6t
Xbit_r108_c86 bl_86 br_86 wl_108 vdd gnd cell_6t
Xbit_r109_c86 bl_86 br_86 wl_109 vdd gnd cell_6t
Xbit_r110_c86 bl_86 br_86 wl_110 vdd gnd cell_6t
Xbit_r111_c86 bl_86 br_86 wl_111 vdd gnd cell_6t
Xbit_r112_c86 bl_86 br_86 wl_112 vdd gnd cell_6t
Xbit_r113_c86 bl_86 br_86 wl_113 vdd gnd cell_6t
Xbit_r114_c86 bl_86 br_86 wl_114 vdd gnd cell_6t
Xbit_r115_c86 bl_86 br_86 wl_115 vdd gnd cell_6t
Xbit_r116_c86 bl_86 br_86 wl_116 vdd gnd cell_6t
Xbit_r117_c86 bl_86 br_86 wl_117 vdd gnd cell_6t
Xbit_r118_c86 bl_86 br_86 wl_118 vdd gnd cell_6t
Xbit_r119_c86 bl_86 br_86 wl_119 vdd gnd cell_6t
Xbit_r120_c86 bl_86 br_86 wl_120 vdd gnd cell_6t
Xbit_r121_c86 bl_86 br_86 wl_121 vdd gnd cell_6t
Xbit_r122_c86 bl_86 br_86 wl_122 vdd gnd cell_6t
Xbit_r123_c86 bl_86 br_86 wl_123 vdd gnd cell_6t
Xbit_r124_c86 bl_86 br_86 wl_124 vdd gnd cell_6t
Xbit_r125_c86 bl_86 br_86 wl_125 vdd gnd cell_6t
Xbit_r126_c86 bl_86 br_86 wl_126 vdd gnd cell_6t
Xbit_r127_c86 bl_86 br_86 wl_127 vdd gnd cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd cell_6t
Xbit_r1_c87 bl_87 br_87 wl_1 vdd gnd cell_6t
Xbit_r2_c87 bl_87 br_87 wl_2 vdd gnd cell_6t
Xbit_r3_c87 bl_87 br_87 wl_3 vdd gnd cell_6t
Xbit_r4_c87 bl_87 br_87 wl_4 vdd gnd cell_6t
Xbit_r5_c87 bl_87 br_87 wl_5 vdd gnd cell_6t
Xbit_r6_c87 bl_87 br_87 wl_6 vdd gnd cell_6t
Xbit_r7_c87 bl_87 br_87 wl_7 vdd gnd cell_6t
Xbit_r8_c87 bl_87 br_87 wl_8 vdd gnd cell_6t
Xbit_r9_c87 bl_87 br_87 wl_9 vdd gnd cell_6t
Xbit_r10_c87 bl_87 br_87 wl_10 vdd gnd cell_6t
Xbit_r11_c87 bl_87 br_87 wl_11 vdd gnd cell_6t
Xbit_r12_c87 bl_87 br_87 wl_12 vdd gnd cell_6t
Xbit_r13_c87 bl_87 br_87 wl_13 vdd gnd cell_6t
Xbit_r14_c87 bl_87 br_87 wl_14 vdd gnd cell_6t
Xbit_r15_c87 bl_87 br_87 wl_15 vdd gnd cell_6t
Xbit_r16_c87 bl_87 br_87 wl_16 vdd gnd cell_6t
Xbit_r17_c87 bl_87 br_87 wl_17 vdd gnd cell_6t
Xbit_r18_c87 bl_87 br_87 wl_18 vdd gnd cell_6t
Xbit_r19_c87 bl_87 br_87 wl_19 vdd gnd cell_6t
Xbit_r20_c87 bl_87 br_87 wl_20 vdd gnd cell_6t
Xbit_r21_c87 bl_87 br_87 wl_21 vdd gnd cell_6t
Xbit_r22_c87 bl_87 br_87 wl_22 vdd gnd cell_6t
Xbit_r23_c87 bl_87 br_87 wl_23 vdd gnd cell_6t
Xbit_r24_c87 bl_87 br_87 wl_24 vdd gnd cell_6t
Xbit_r25_c87 bl_87 br_87 wl_25 vdd gnd cell_6t
Xbit_r26_c87 bl_87 br_87 wl_26 vdd gnd cell_6t
Xbit_r27_c87 bl_87 br_87 wl_27 vdd gnd cell_6t
Xbit_r28_c87 bl_87 br_87 wl_28 vdd gnd cell_6t
Xbit_r29_c87 bl_87 br_87 wl_29 vdd gnd cell_6t
Xbit_r30_c87 bl_87 br_87 wl_30 vdd gnd cell_6t
Xbit_r31_c87 bl_87 br_87 wl_31 vdd gnd cell_6t
Xbit_r32_c87 bl_87 br_87 wl_32 vdd gnd cell_6t
Xbit_r33_c87 bl_87 br_87 wl_33 vdd gnd cell_6t
Xbit_r34_c87 bl_87 br_87 wl_34 vdd gnd cell_6t
Xbit_r35_c87 bl_87 br_87 wl_35 vdd gnd cell_6t
Xbit_r36_c87 bl_87 br_87 wl_36 vdd gnd cell_6t
Xbit_r37_c87 bl_87 br_87 wl_37 vdd gnd cell_6t
Xbit_r38_c87 bl_87 br_87 wl_38 vdd gnd cell_6t
Xbit_r39_c87 bl_87 br_87 wl_39 vdd gnd cell_6t
Xbit_r40_c87 bl_87 br_87 wl_40 vdd gnd cell_6t
Xbit_r41_c87 bl_87 br_87 wl_41 vdd gnd cell_6t
Xbit_r42_c87 bl_87 br_87 wl_42 vdd gnd cell_6t
Xbit_r43_c87 bl_87 br_87 wl_43 vdd gnd cell_6t
Xbit_r44_c87 bl_87 br_87 wl_44 vdd gnd cell_6t
Xbit_r45_c87 bl_87 br_87 wl_45 vdd gnd cell_6t
Xbit_r46_c87 bl_87 br_87 wl_46 vdd gnd cell_6t
Xbit_r47_c87 bl_87 br_87 wl_47 vdd gnd cell_6t
Xbit_r48_c87 bl_87 br_87 wl_48 vdd gnd cell_6t
Xbit_r49_c87 bl_87 br_87 wl_49 vdd gnd cell_6t
Xbit_r50_c87 bl_87 br_87 wl_50 vdd gnd cell_6t
Xbit_r51_c87 bl_87 br_87 wl_51 vdd gnd cell_6t
Xbit_r52_c87 bl_87 br_87 wl_52 vdd gnd cell_6t
Xbit_r53_c87 bl_87 br_87 wl_53 vdd gnd cell_6t
Xbit_r54_c87 bl_87 br_87 wl_54 vdd gnd cell_6t
Xbit_r55_c87 bl_87 br_87 wl_55 vdd gnd cell_6t
Xbit_r56_c87 bl_87 br_87 wl_56 vdd gnd cell_6t
Xbit_r57_c87 bl_87 br_87 wl_57 vdd gnd cell_6t
Xbit_r58_c87 bl_87 br_87 wl_58 vdd gnd cell_6t
Xbit_r59_c87 bl_87 br_87 wl_59 vdd gnd cell_6t
Xbit_r60_c87 bl_87 br_87 wl_60 vdd gnd cell_6t
Xbit_r61_c87 bl_87 br_87 wl_61 vdd gnd cell_6t
Xbit_r62_c87 bl_87 br_87 wl_62 vdd gnd cell_6t
Xbit_r63_c87 bl_87 br_87 wl_63 vdd gnd cell_6t
Xbit_r64_c87 bl_87 br_87 wl_64 vdd gnd cell_6t
Xbit_r65_c87 bl_87 br_87 wl_65 vdd gnd cell_6t
Xbit_r66_c87 bl_87 br_87 wl_66 vdd gnd cell_6t
Xbit_r67_c87 bl_87 br_87 wl_67 vdd gnd cell_6t
Xbit_r68_c87 bl_87 br_87 wl_68 vdd gnd cell_6t
Xbit_r69_c87 bl_87 br_87 wl_69 vdd gnd cell_6t
Xbit_r70_c87 bl_87 br_87 wl_70 vdd gnd cell_6t
Xbit_r71_c87 bl_87 br_87 wl_71 vdd gnd cell_6t
Xbit_r72_c87 bl_87 br_87 wl_72 vdd gnd cell_6t
Xbit_r73_c87 bl_87 br_87 wl_73 vdd gnd cell_6t
Xbit_r74_c87 bl_87 br_87 wl_74 vdd gnd cell_6t
Xbit_r75_c87 bl_87 br_87 wl_75 vdd gnd cell_6t
Xbit_r76_c87 bl_87 br_87 wl_76 vdd gnd cell_6t
Xbit_r77_c87 bl_87 br_87 wl_77 vdd gnd cell_6t
Xbit_r78_c87 bl_87 br_87 wl_78 vdd gnd cell_6t
Xbit_r79_c87 bl_87 br_87 wl_79 vdd gnd cell_6t
Xbit_r80_c87 bl_87 br_87 wl_80 vdd gnd cell_6t
Xbit_r81_c87 bl_87 br_87 wl_81 vdd gnd cell_6t
Xbit_r82_c87 bl_87 br_87 wl_82 vdd gnd cell_6t
Xbit_r83_c87 bl_87 br_87 wl_83 vdd gnd cell_6t
Xbit_r84_c87 bl_87 br_87 wl_84 vdd gnd cell_6t
Xbit_r85_c87 bl_87 br_87 wl_85 vdd gnd cell_6t
Xbit_r86_c87 bl_87 br_87 wl_86 vdd gnd cell_6t
Xbit_r87_c87 bl_87 br_87 wl_87 vdd gnd cell_6t
Xbit_r88_c87 bl_87 br_87 wl_88 vdd gnd cell_6t
Xbit_r89_c87 bl_87 br_87 wl_89 vdd gnd cell_6t
Xbit_r90_c87 bl_87 br_87 wl_90 vdd gnd cell_6t
Xbit_r91_c87 bl_87 br_87 wl_91 vdd gnd cell_6t
Xbit_r92_c87 bl_87 br_87 wl_92 vdd gnd cell_6t
Xbit_r93_c87 bl_87 br_87 wl_93 vdd gnd cell_6t
Xbit_r94_c87 bl_87 br_87 wl_94 vdd gnd cell_6t
Xbit_r95_c87 bl_87 br_87 wl_95 vdd gnd cell_6t
Xbit_r96_c87 bl_87 br_87 wl_96 vdd gnd cell_6t
Xbit_r97_c87 bl_87 br_87 wl_97 vdd gnd cell_6t
Xbit_r98_c87 bl_87 br_87 wl_98 vdd gnd cell_6t
Xbit_r99_c87 bl_87 br_87 wl_99 vdd gnd cell_6t
Xbit_r100_c87 bl_87 br_87 wl_100 vdd gnd cell_6t
Xbit_r101_c87 bl_87 br_87 wl_101 vdd gnd cell_6t
Xbit_r102_c87 bl_87 br_87 wl_102 vdd gnd cell_6t
Xbit_r103_c87 bl_87 br_87 wl_103 vdd gnd cell_6t
Xbit_r104_c87 bl_87 br_87 wl_104 vdd gnd cell_6t
Xbit_r105_c87 bl_87 br_87 wl_105 vdd gnd cell_6t
Xbit_r106_c87 bl_87 br_87 wl_106 vdd gnd cell_6t
Xbit_r107_c87 bl_87 br_87 wl_107 vdd gnd cell_6t
Xbit_r108_c87 bl_87 br_87 wl_108 vdd gnd cell_6t
Xbit_r109_c87 bl_87 br_87 wl_109 vdd gnd cell_6t
Xbit_r110_c87 bl_87 br_87 wl_110 vdd gnd cell_6t
Xbit_r111_c87 bl_87 br_87 wl_111 vdd gnd cell_6t
Xbit_r112_c87 bl_87 br_87 wl_112 vdd gnd cell_6t
Xbit_r113_c87 bl_87 br_87 wl_113 vdd gnd cell_6t
Xbit_r114_c87 bl_87 br_87 wl_114 vdd gnd cell_6t
Xbit_r115_c87 bl_87 br_87 wl_115 vdd gnd cell_6t
Xbit_r116_c87 bl_87 br_87 wl_116 vdd gnd cell_6t
Xbit_r117_c87 bl_87 br_87 wl_117 vdd gnd cell_6t
Xbit_r118_c87 bl_87 br_87 wl_118 vdd gnd cell_6t
Xbit_r119_c87 bl_87 br_87 wl_119 vdd gnd cell_6t
Xbit_r120_c87 bl_87 br_87 wl_120 vdd gnd cell_6t
Xbit_r121_c87 bl_87 br_87 wl_121 vdd gnd cell_6t
Xbit_r122_c87 bl_87 br_87 wl_122 vdd gnd cell_6t
Xbit_r123_c87 bl_87 br_87 wl_123 vdd gnd cell_6t
Xbit_r124_c87 bl_87 br_87 wl_124 vdd gnd cell_6t
Xbit_r125_c87 bl_87 br_87 wl_125 vdd gnd cell_6t
Xbit_r126_c87 bl_87 br_87 wl_126 vdd gnd cell_6t
Xbit_r127_c87 bl_87 br_87 wl_127 vdd gnd cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd cell_6t
Xbit_r1_c88 bl_88 br_88 wl_1 vdd gnd cell_6t
Xbit_r2_c88 bl_88 br_88 wl_2 vdd gnd cell_6t
Xbit_r3_c88 bl_88 br_88 wl_3 vdd gnd cell_6t
Xbit_r4_c88 bl_88 br_88 wl_4 vdd gnd cell_6t
Xbit_r5_c88 bl_88 br_88 wl_5 vdd gnd cell_6t
Xbit_r6_c88 bl_88 br_88 wl_6 vdd gnd cell_6t
Xbit_r7_c88 bl_88 br_88 wl_7 vdd gnd cell_6t
Xbit_r8_c88 bl_88 br_88 wl_8 vdd gnd cell_6t
Xbit_r9_c88 bl_88 br_88 wl_9 vdd gnd cell_6t
Xbit_r10_c88 bl_88 br_88 wl_10 vdd gnd cell_6t
Xbit_r11_c88 bl_88 br_88 wl_11 vdd gnd cell_6t
Xbit_r12_c88 bl_88 br_88 wl_12 vdd gnd cell_6t
Xbit_r13_c88 bl_88 br_88 wl_13 vdd gnd cell_6t
Xbit_r14_c88 bl_88 br_88 wl_14 vdd gnd cell_6t
Xbit_r15_c88 bl_88 br_88 wl_15 vdd gnd cell_6t
Xbit_r16_c88 bl_88 br_88 wl_16 vdd gnd cell_6t
Xbit_r17_c88 bl_88 br_88 wl_17 vdd gnd cell_6t
Xbit_r18_c88 bl_88 br_88 wl_18 vdd gnd cell_6t
Xbit_r19_c88 bl_88 br_88 wl_19 vdd gnd cell_6t
Xbit_r20_c88 bl_88 br_88 wl_20 vdd gnd cell_6t
Xbit_r21_c88 bl_88 br_88 wl_21 vdd gnd cell_6t
Xbit_r22_c88 bl_88 br_88 wl_22 vdd gnd cell_6t
Xbit_r23_c88 bl_88 br_88 wl_23 vdd gnd cell_6t
Xbit_r24_c88 bl_88 br_88 wl_24 vdd gnd cell_6t
Xbit_r25_c88 bl_88 br_88 wl_25 vdd gnd cell_6t
Xbit_r26_c88 bl_88 br_88 wl_26 vdd gnd cell_6t
Xbit_r27_c88 bl_88 br_88 wl_27 vdd gnd cell_6t
Xbit_r28_c88 bl_88 br_88 wl_28 vdd gnd cell_6t
Xbit_r29_c88 bl_88 br_88 wl_29 vdd gnd cell_6t
Xbit_r30_c88 bl_88 br_88 wl_30 vdd gnd cell_6t
Xbit_r31_c88 bl_88 br_88 wl_31 vdd gnd cell_6t
Xbit_r32_c88 bl_88 br_88 wl_32 vdd gnd cell_6t
Xbit_r33_c88 bl_88 br_88 wl_33 vdd gnd cell_6t
Xbit_r34_c88 bl_88 br_88 wl_34 vdd gnd cell_6t
Xbit_r35_c88 bl_88 br_88 wl_35 vdd gnd cell_6t
Xbit_r36_c88 bl_88 br_88 wl_36 vdd gnd cell_6t
Xbit_r37_c88 bl_88 br_88 wl_37 vdd gnd cell_6t
Xbit_r38_c88 bl_88 br_88 wl_38 vdd gnd cell_6t
Xbit_r39_c88 bl_88 br_88 wl_39 vdd gnd cell_6t
Xbit_r40_c88 bl_88 br_88 wl_40 vdd gnd cell_6t
Xbit_r41_c88 bl_88 br_88 wl_41 vdd gnd cell_6t
Xbit_r42_c88 bl_88 br_88 wl_42 vdd gnd cell_6t
Xbit_r43_c88 bl_88 br_88 wl_43 vdd gnd cell_6t
Xbit_r44_c88 bl_88 br_88 wl_44 vdd gnd cell_6t
Xbit_r45_c88 bl_88 br_88 wl_45 vdd gnd cell_6t
Xbit_r46_c88 bl_88 br_88 wl_46 vdd gnd cell_6t
Xbit_r47_c88 bl_88 br_88 wl_47 vdd gnd cell_6t
Xbit_r48_c88 bl_88 br_88 wl_48 vdd gnd cell_6t
Xbit_r49_c88 bl_88 br_88 wl_49 vdd gnd cell_6t
Xbit_r50_c88 bl_88 br_88 wl_50 vdd gnd cell_6t
Xbit_r51_c88 bl_88 br_88 wl_51 vdd gnd cell_6t
Xbit_r52_c88 bl_88 br_88 wl_52 vdd gnd cell_6t
Xbit_r53_c88 bl_88 br_88 wl_53 vdd gnd cell_6t
Xbit_r54_c88 bl_88 br_88 wl_54 vdd gnd cell_6t
Xbit_r55_c88 bl_88 br_88 wl_55 vdd gnd cell_6t
Xbit_r56_c88 bl_88 br_88 wl_56 vdd gnd cell_6t
Xbit_r57_c88 bl_88 br_88 wl_57 vdd gnd cell_6t
Xbit_r58_c88 bl_88 br_88 wl_58 vdd gnd cell_6t
Xbit_r59_c88 bl_88 br_88 wl_59 vdd gnd cell_6t
Xbit_r60_c88 bl_88 br_88 wl_60 vdd gnd cell_6t
Xbit_r61_c88 bl_88 br_88 wl_61 vdd gnd cell_6t
Xbit_r62_c88 bl_88 br_88 wl_62 vdd gnd cell_6t
Xbit_r63_c88 bl_88 br_88 wl_63 vdd gnd cell_6t
Xbit_r64_c88 bl_88 br_88 wl_64 vdd gnd cell_6t
Xbit_r65_c88 bl_88 br_88 wl_65 vdd gnd cell_6t
Xbit_r66_c88 bl_88 br_88 wl_66 vdd gnd cell_6t
Xbit_r67_c88 bl_88 br_88 wl_67 vdd gnd cell_6t
Xbit_r68_c88 bl_88 br_88 wl_68 vdd gnd cell_6t
Xbit_r69_c88 bl_88 br_88 wl_69 vdd gnd cell_6t
Xbit_r70_c88 bl_88 br_88 wl_70 vdd gnd cell_6t
Xbit_r71_c88 bl_88 br_88 wl_71 vdd gnd cell_6t
Xbit_r72_c88 bl_88 br_88 wl_72 vdd gnd cell_6t
Xbit_r73_c88 bl_88 br_88 wl_73 vdd gnd cell_6t
Xbit_r74_c88 bl_88 br_88 wl_74 vdd gnd cell_6t
Xbit_r75_c88 bl_88 br_88 wl_75 vdd gnd cell_6t
Xbit_r76_c88 bl_88 br_88 wl_76 vdd gnd cell_6t
Xbit_r77_c88 bl_88 br_88 wl_77 vdd gnd cell_6t
Xbit_r78_c88 bl_88 br_88 wl_78 vdd gnd cell_6t
Xbit_r79_c88 bl_88 br_88 wl_79 vdd gnd cell_6t
Xbit_r80_c88 bl_88 br_88 wl_80 vdd gnd cell_6t
Xbit_r81_c88 bl_88 br_88 wl_81 vdd gnd cell_6t
Xbit_r82_c88 bl_88 br_88 wl_82 vdd gnd cell_6t
Xbit_r83_c88 bl_88 br_88 wl_83 vdd gnd cell_6t
Xbit_r84_c88 bl_88 br_88 wl_84 vdd gnd cell_6t
Xbit_r85_c88 bl_88 br_88 wl_85 vdd gnd cell_6t
Xbit_r86_c88 bl_88 br_88 wl_86 vdd gnd cell_6t
Xbit_r87_c88 bl_88 br_88 wl_87 vdd gnd cell_6t
Xbit_r88_c88 bl_88 br_88 wl_88 vdd gnd cell_6t
Xbit_r89_c88 bl_88 br_88 wl_89 vdd gnd cell_6t
Xbit_r90_c88 bl_88 br_88 wl_90 vdd gnd cell_6t
Xbit_r91_c88 bl_88 br_88 wl_91 vdd gnd cell_6t
Xbit_r92_c88 bl_88 br_88 wl_92 vdd gnd cell_6t
Xbit_r93_c88 bl_88 br_88 wl_93 vdd gnd cell_6t
Xbit_r94_c88 bl_88 br_88 wl_94 vdd gnd cell_6t
Xbit_r95_c88 bl_88 br_88 wl_95 vdd gnd cell_6t
Xbit_r96_c88 bl_88 br_88 wl_96 vdd gnd cell_6t
Xbit_r97_c88 bl_88 br_88 wl_97 vdd gnd cell_6t
Xbit_r98_c88 bl_88 br_88 wl_98 vdd gnd cell_6t
Xbit_r99_c88 bl_88 br_88 wl_99 vdd gnd cell_6t
Xbit_r100_c88 bl_88 br_88 wl_100 vdd gnd cell_6t
Xbit_r101_c88 bl_88 br_88 wl_101 vdd gnd cell_6t
Xbit_r102_c88 bl_88 br_88 wl_102 vdd gnd cell_6t
Xbit_r103_c88 bl_88 br_88 wl_103 vdd gnd cell_6t
Xbit_r104_c88 bl_88 br_88 wl_104 vdd gnd cell_6t
Xbit_r105_c88 bl_88 br_88 wl_105 vdd gnd cell_6t
Xbit_r106_c88 bl_88 br_88 wl_106 vdd gnd cell_6t
Xbit_r107_c88 bl_88 br_88 wl_107 vdd gnd cell_6t
Xbit_r108_c88 bl_88 br_88 wl_108 vdd gnd cell_6t
Xbit_r109_c88 bl_88 br_88 wl_109 vdd gnd cell_6t
Xbit_r110_c88 bl_88 br_88 wl_110 vdd gnd cell_6t
Xbit_r111_c88 bl_88 br_88 wl_111 vdd gnd cell_6t
Xbit_r112_c88 bl_88 br_88 wl_112 vdd gnd cell_6t
Xbit_r113_c88 bl_88 br_88 wl_113 vdd gnd cell_6t
Xbit_r114_c88 bl_88 br_88 wl_114 vdd gnd cell_6t
Xbit_r115_c88 bl_88 br_88 wl_115 vdd gnd cell_6t
Xbit_r116_c88 bl_88 br_88 wl_116 vdd gnd cell_6t
Xbit_r117_c88 bl_88 br_88 wl_117 vdd gnd cell_6t
Xbit_r118_c88 bl_88 br_88 wl_118 vdd gnd cell_6t
Xbit_r119_c88 bl_88 br_88 wl_119 vdd gnd cell_6t
Xbit_r120_c88 bl_88 br_88 wl_120 vdd gnd cell_6t
Xbit_r121_c88 bl_88 br_88 wl_121 vdd gnd cell_6t
Xbit_r122_c88 bl_88 br_88 wl_122 vdd gnd cell_6t
Xbit_r123_c88 bl_88 br_88 wl_123 vdd gnd cell_6t
Xbit_r124_c88 bl_88 br_88 wl_124 vdd gnd cell_6t
Xbit_r125_c88 bl_88 br_88 wl_125 vdd gnd cell_6t
Xbit_r126_c88 bl_88 br_88 wl_126 vdd gnd cell_6t
Xbit_r127_c88 bl_88 br_88 wl_127 vdd gnd cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd cell_6t
Xbit_r1_c89 bl_89 br_89 wl_1 vdd gnd cell_6t
Xbit_r2_c89 bl_89 br_89 wl_2 vdd gnd cell_6t
Xbit_r3_c89 bl_89 br_89 wl_3 vdd gnd cell_6t
Xbit_r4_c89 bl_89 br_89 wl_4 vdd gnd cell_6t
Xbit_r5_c89 bl_89 br_89 wl_5 vdd gnd cell_6t
Xbit_r6_c89 bl_89 br_89 wl_6 vdd gnd cell_6t
Xbit_r7_c89 bl_89 br_89 wl_7 vdd gnd cell_6t
Xbit_r8_c89 bl_89 br_89 wl_8 vdd gnd cell_6t
Xbit_r9_c89 bl_89 br_89 wl_9 vdd gnd cell_6t
Xbit_r10_c89 bl_89 br_89 wl_10 vdd gnd cell_6t
Xbit_r11_c89 bl_89 br_89 wl_11 vdd gnd cell_6t
Xbit_r12_c89 bl_89 br_89 wl_12 vdd gnd cell_6t
Xbit_r13_c89 bl_89 br_89 wl_13 vdd gnd cell_6t
Xbit_r14_c89 bl_89 br_89 wl_14 vdd gnd cell_6t
Xbit_r15_c89 bl_89 br_89 wl_15 vdd gnd cell_6t
Xbit_r16_c89 bl_89 br_89 wl_16 vdd gnd cell_6t
Xbit_r17_c89 bl_89 br_89 wl_17 vdd gnd cell_6t
Xbit_r18_c89 bl_89 br_89 wl_18 vdd gnd cell_6t
Xbit_r19_c89 bl_89 br_89 wl_19 vdd gnd cell_6t
Xbit_r20_c89 bl_89 br_89 wl_20 vdd gnd cell_6t
Xbit_r21_c89 bl_89 br_89 wl_21 vdd gnd cell_6t
Xbit_r22_c89 bl_89 br_89 wl_22 vdd gnd cell_6t
Xbit_r23_c89 bl_89 br_89 wl_23 vdd gnd cell_6t
Xbit_r24_c89 bl_89 br_89 wl_24 vdd gnd cell_6t
Xbit_r25_c89 bl_89 br_89 wl_25 vdd gnd cell_6t
Xbit_r26_c89 bl_89 br_89 wl_26 vdd gnd cell_6t
Xbit_r27_c89 bl_89 br_89 wl_27 vdd gnd cell_6t
Xbit_r28_c89 bl_89 br_89 wl_28 vdd gnd cell_6t
Xbit_r29_c89 bl_89 br_89 wl_29 vdd gnd cell_6t
Xbit_r30_c89 bl_89 br_89 wl_30 vdd gnd cell_6t
Xbit_r31_c89 bl_89 br_89 wl_31 vdd gnd cell_6t
Xbit_r32_c89 bl_89 br_89 wl_32 vdd gnd cell_6t
Xbit_r33_c89 bl_89 br_89 wl_33 vdd gnd cell_6t
Xbit_r34_c89 bl_89 br_89 wl_34 vdd gnd cell_6t
Xbit_r35_c89 bl_89 br_89 wl_35 vdd gnd cell_6t
Xbit_r36_c89 bl_89 br_89 wl_36 vdd gnd cell_6t
Xbit_r37_c89 bl_89 br_89 wl_37 vdd gnd cell_6t
Xbit_r38_c89 bl_89 br_89 wl_38 vdd gnd cell_6t
Xbit_r39_c89 bl_89 br_89 wl_39 vdd gnd cell_6t
Xbit_r40_c89 bl_89 br_89 wl_40 vdd gnd cell_6t
Xbit_r41_c89 bl_89 br_89 wl_41 vdd gnd cell_6t
Xbit_r42_c89 bl_89 br_89 wl_42 vdd gnd cell_6t
Xbit_r43_c89 bl_89 br_89 wl_43 vdd gnd cell_6t
Xbit_r44_c89 bl_89 br_89 wl_44 vdd gnd cell_6t
Xbit_r45_c89 bl_89 br_89 wl_45 vdd gnd cell_6t
Xbit_r46_c89 bl_89 br_89 wl_46 vdd gnd cell_6t
Xbit_r47_c89 bl_89 br_89 wl_47 vdd gnd cell_6t
Xbit_r48_c89 bl_89 br_89 wl_48 vdd gnd cell_6t
Xbit_r49_c89 bl_89 br_89 wl_49 vdd gnd cell_6t
Xbit_r50_c89 bl_89 br_89 wl_50 vdd gnd cell_6t
Xbit_r51_c89 bl_89 br_89 wl_51 vdd gnd cell_6t
Xbit_r52_c89 bl_89 br_89 wl_52 vdd gnd cell_6t
Xbit_r53_c89 bl_89 br_89 wl_53 vdd gnd cell_6t
Xbit_r54_c89 bl_89 br_89 wl_54 vdd gnd cell_6t
Xbit_r55_c89 bl_89 br_89 wl_55 vdd gnd cell_6t
Xbit_r56_c89 bl_89 br_89 wl_56 vdd gnd cell_6t
Xbit_r57_c89 bl_89 br_89 wl_57 vdd gnd cell_6t
Xbit_r58_c89 bl_89 br_89 wl_58 vdd gnd cell_6t
Xbit_r59_c89 bl_89 br_89 wl_59 vdd gnd cell_6t
Xbit_r60_c89 bl_89 br_89 wl_60 vdd gnd cell_6t
Xbit_r61_c89 bl_89 br_89 wl_61 vdd gnd cell_6t
Xbit_r62_c89 bl_89 br_89 wl_62 vdd gnd cell_6t
Xbit_r63_c89 bl_89 br_89 wl_63 vdd gnd cell_6t
Xbit_r64_c89 bl_89 br_89 wl_64 vdd gnd cell_6t
Xbit_r65_c89 bl_89 br_89 wl_65 vdd gnd cell_6t
Xbit_r66_c89 bl_89 br_89 wl_66 vdd gnd cell_6t
Xbit_r67_c89 bl_89 br_89 wl_67 vdd gnd cell_6t
Xbit_r68_c89 bl_89 br_89 wl_68 vdd gnd cell_6t
Xbit_r69_c89 bl_89 br_89 wl_69 vdd gnd cell_6t
Xbit_r70_c89 bl_89 br_89 wl_70 vdd gnd cell_6t
Xbit_r71_c89 bl_89 br_89 wl_71 vdd gnd cell_6t
Xbit_r72_c89 bl_89 br_89 wl_72 vdd gnd cell_6t
Xbit_r73_c89 bl_89 br_89 wl_73 vdd gnd cell_6t
Xbit_r74_c89 bl_89 br_89 wl_74 vdd gnd cell_6t
Xbit_r75_c89 bl_89 br_89 wl_75 vdd gnd cell_6t
Xbit_r76_c89 bl_89 br_89 wl_76 vdd gnd cell_6t
Xbit_r77_c89 bl_89 br_89 wl_77 vdd gnd cell_6t
Xbit_r78_c89 bl_89 br_89 wl_78 vdd gnd cell_6t
Xbit_r79_c89 bl_89 br_89 wl_79 vdd gnd cell_6t
Xbit_r80_c89 bl_89 br_89 wl_80 vdd gnd cell_6t
Xbit_r81_c89 bl_89 br_89 wl_81 vdd gnd cell_6t
Xbit_r82_c89 bl_89 br_89 wl_82 vdd gnd cell_6t
Xbit_r83_c89 bl_89 br_89 wl_83 vdd gnd cell_6t
Xbit_r84_c89 bl_89 br_89 wl_84 vdd gnd cell_6t
Xbit_r85_c89 bl_89 br_89 wl_85 vdd gnd cell_6t
Xbit_r86_c89 bl_89 br_89 wl_86 vdd gnd cell_6t
Xbit_r87_c89 bl_89 br_89 wl_87 vdd gnd cell_6t
Xbit_r88_c89 bl_89 br_89 wl_88 vdd gnd cell_6t
Xbit_r89_c89 bl_89 br_89 wl_89 vdd gnd cell_6t
Xbit_r90_c89 bl_89 br_89 wl_90 vdd gnd cell_6t
Xbit_r91_c89 bl_89 br_89 wl_91 vdd gnd cell_6t
Xbit_r92_c89 bl_89 br_89 wl_92 vdd gnd cell_6t
Xbit_r93_c89 bl_89 br_89 wl_93 vdd gnd cell_6t
Xbit_r94_c89 bl_89 br_89 wl_94 vdd gnd cell_6t
Xbit_r95_c89 bl_89 br_89 wl_95 vdd gnd cell_6t
Xbit_r96_c89 bl_89 br_89 wl_96 vdd gnd cell_6t
Xbit_r97_c89 bl_89 br_89 wl_97 vdd gnd cell_6t
Xbit_r98_c89 bl_89 br_89 wl_98 vdd gnd cell_6t
Xbit_r99_c89 bl_89 br_89 wl_99 vdd gnd cell_6t
Xbit_r100_c89 bl_89 br_89 wl_100 vdd gnd cell_6t
Xbit_r101_c89 bl_89 br_89 wl_101 vdd gnd cell_6t
Xbit_r102_c89 bl_89 br_89 wl_102 vdd gnd cell_6t
Xbit_r103_c89 bl_89 br_89 wl_103 vdd gnd cell_6t
Xbit_r104_c89 bl_89 br_89 wl_104 vdd gnd cell_6t
Xbit_r105_c89 bl_89 br_89 wl_105 vdd gnd cell_6t
Xbit_r106_c89 bl_89 br_89 wl_106 vdd gnd cell_6t
Xbit_r107_c89 bl_89 br_89 wl_107 vdd gnd cell_6t
Xbit_r108_c89 bl_89 br_89 wl_108 vdd gnd cell_6t
Xbit_r109_c89 bl_89 br_89 wl_109 vdd gnd cell_6t
Xbit_r110_c89 bl_89 br_89 wl_110 vdd gnd cell_6t
Xbit_r111_c89 bl_89 br_89 wl_111 vdd gnd cell_6t
Xbit_r112_c89 bl_89 br_89 wl_112 vdd gnd cell_6t
Xbit_r113_c89 bl_89 br_89 wl_113 vdd gnd cell_6t
Xbit_r114_c89 bl_89 br_89 wl_114 vdd gnd cell_6t
Xbit_r115_c89 bl_89 br_89 wl_115 vdd gnd cell_6t
Xbit_r116_c89 bl_89 br_89 wl_116 vdd gnd cell_6t
Xbit_r117_c89 bl_89 br_89 wl_117 vdd gnd cell_6t
Xbit_r118_c89 bl_89 br_89 wl_118 vdd gnd cell_6t
Xbit_r119_c89 bl_89 br_89 wl_119 vdd gnd cell_6t
Xbit_r120_c89 bl_89 br_89 wl_120 vdd gnd cell_6t
Xbit_r121_c89 bl_89 br_89 wl_121 vdd gnd cell_6t
Xbit_r122_c89 bl_89 br_89 wl_122 vdd gnd cell_6t
Xbit_r123_c89 bl_89 br_89 wl_123 vdd gnd cell_6t
Xbit_r124_c89 bl_89 br_89 wl_124 vdd gnd cell_6t
Xbit_r125_c89 bl_89 br_89 wl_125 vdd gnd cell_6t
Xbit_r126_c89 bl_89 br_89 wl_126 vdd gnd cell_6t
Xbit_r127_c89 bl_89 br_89 wl_127 vdd gnd cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd cell_6t
Xbit_r1_c90 bl_90 br_90 wl_1 vdd gnd cell_6t
Xbit_r2_c90 bl_90 br_90 wl_2 vdd gnd cell_6t
Xbit_r3_c90 bl_90 br_90 wl_3 vdd gnd cell_6t
Xbit_r4_c90 bl_90 br_90 wl_4 vdd gnd cell_6t
Xbit_r5_c90 bl_90 br_90 wl_5 vdd gnd cell_6t
Xbit_r6_c90 bl_90 br_90 wl_6 vdd gnd cell_6t
Xbit_r7_c90 bl_90 br_90 wl_7 vdd gnd cell_6t
Xbit_r8_c90 bl_90 br_90 wl_8 vdd gnd cell_6t
Xbit_r9_c90 bl_90 br_90 wl_9 vdd gnd cell_6t
Xbit_r10_c90 bl_90 br_90 wl_10 vdd gnd cell_6t
Xbit_r11_c90 bl_90 br_90 wl_11 vdd gnd cell_6t
Xbit_r12_c90 bl_90 br_90 wl_12 vdd gnd cell_6t
Xbit_r13_c90 bl_90 br_90 wl_13 vdd gnd cell_6t
Xbit_r14_c90 bl_90 br_90 wl_14 vdd gnd cell_6t
Xbit_r15_c90 bl_90 br_90 wl_15 vdd gnd cell_6t
Xbit_r16_c90 bl_90 br_90 wl_16 vdd gnd cell_6t
Xbit_r17_c90 bl_90 br_90 wl_17 vdd gnd cell_6t
Xbit_r18_c90 bl_90 br_90 wl_18 vdd gnd cell_6t
Xbit_r19_c90 bl_90 br_90 wl_19 vdd gnd cell_6t
Xbit_r20_c90 bl_90 br_90 wl_20 vdd gnd cell_6t
Xbit_r21_c90 bl_90 br_90 wl_21 vdd gnd cell_6t
Xbit_r22_c90 bl_90 br_90 wl_22 vdd gnd cell_6t
Xbit_r23_c90 bl_90 br_90 wl_23 vdd gnd cell_6t
Xbit_r24_c90 bl_90 br_90 wl_24 vdd gnd cell_6t
Xbit_r25_c90 bl_90 br_90 wl_25 vdd gnd cell_6t
Xbit_r26_c90 bl_90 br_90 wl_26 vdd gnd cell_6t
Xbit_r27_c90 bl_90 br_90 wl_27 vdd gnd cell_6t
Xbit_r28_c90 bl_90 br_90 wl_28 vdd gnd cell_6t
Xbit_r29_c90 bl_90 br_90 wl_29 vdd gnd cell_6t
Xbit_r30_c90 bl_90 br_90 wl_30 vdd gnd cell_6t
Xbit_r31_c90 bl_90 br_90 wl_31 vdd gnd cell_6t
Xbit_r32_c90 bl_90 br_90 wl_32 vdd gnd cell_6t
Xbit_r33_c90 bl_90 br_90 wl_33 vdd gnd cell_6t
Xbit_r34_c90 bl_90 br_90 wl_34 vdd gnd cell_6t
Xbit_r35_c90 bl_90 br_90 wl_35 vdd gnd cell_6t
Xbit_r36_c90 bl_90 br_90 wl_36 vdd gnd cell_6t
Xbit_r37_c90 bl_90 br_90 wl_37 vdd gnd cell_6t
Xbit_r38_c90 bl_90 br_90 wl_38 vdd gnd cell_6t
Xbit_r39_c90 bl_90 br_90 wl_39 vdd gnd cell_6t
Xbit_r40_c90 bl_90 br_90 wl_40 vdd gnd cell_6t
Xbit_r41_c90 bl_90 br_90 wl_41 vdd gnd cell_6t
Xbit_r42_c90 bl_90 br_90 wl_42 vdd gnd cell_6t
Xbit_r43_c90 bl_90 br_90 wl_43 vdd gnd cell_6t
Xbit_r44_c90 bl_90 br_90 wl_44 vdd gnd cell_6t
Xbit_r45_c90 bl_90 br_90 wl_45 vdd gnd cell_6t
Xbit_r46_c90 bl_90 br_90 wl_46 vdd gnd cell_6t
Xbit_r47_c90 bl_90 br_90 wl_47 vdd gnd cell_6t
Xbit_r48_c90 bl_90 br_90 wl_48 vdd gnd cell_6t
Xbit_r49_c90 bl_90 br_90 wl_49 vdd gnd cell_6t
Xbit_r50_c90 bl_90 br_90 wl_50 vdd gnd cell_6t
Xbit_r51_c90 bl_90 br_90 wl_51 vdd gnd cell_6t
Xbit_r52_c90 bl_90 br_90 wl_52 vdd gnd cell_6t
Xbit_r53_c90 bl_90 br_90 wl_53 vdd gnd cell_6t
Xbit_r54_c90 bl_90 br_90 wl_54 vdd gnd cell_6t
Xbit_r55_c90 bl_90 br_90 wl_55 vdd gnd cell_6t
Xbit_r56_c90 bl_90 br_90 wl_56 vdd gnd cell_6t
Xbit_r57_c90 bl_90 br_90 wl_57 vdd gnd cell_6t
Xbit_r58_c90 bl_90 br_90 wl_58 vdd gnd cell_6t
Xbit_r59_c90 bl_90 br_90 wl_59 vdd gnd cell_6t
Xbit_r60_c90 bl_90 br_90 wl_60 vdd gnd cell_6t
Xbit_r61_c90 bl_90 br_90 wl_61 vdd gnd cell_6t
Xbit_r62_c90 bl_90 br_90 wl_62 vdd gnd cell_6t
Xbit_r63_c90 bl_90 br_90 wl_63 vdd gnd cell_6t
Xbit_r64_c90 bl_90 br_90 wl_64 vdd gnd cell_6t
Xbit_r65_c90 bl_90 br_90 wl_65 vdd gnd cell_6t
Xbit_r66_c90 bl_90 br_90 wl_66 vdd gnd cell_6t
Xbit_r67_c90 bl_90 br_90 wl_67 vdd gnd cell_6t
Xbit_r68_c90 bl_90 br_90 wl_68 vdd gnd cell_6t
Xbit_r69_c90 bl_90 br_90 wl_69 vdd gnd cell_6t
Xbit_r70_c90 bl_90 br_90 wl_70 vdd gnd cell_6t
Xbit_r71_c90 bl_90 br_90 wl_71 vdd gnd cell_6t
Xbit_r72_c90 bl_90 br_90 wl_72 vdd gnd cell_6t
Xbit_r73_c90 bl_90 br_90 wl_73 vdd gnd cell_6t
Xbit_r74_c90 bl_90 br_90 wl_74 vdd gnd cell_6t
Xbit_r75_c90 bl_90 br_90 wl_75 vdd gnd cell_6t
Xbit_r76_c90 bl_90 br_90 wl_76 vdd gnd cell_6t
Xbit_r77_c90 bl_90 br_90 wl_77 vdd gnd cell_6t
Xbit_r78_c90 bl_90 br_90 wl_78 vdd gnd cell_6t
Xbit_r79_c90 bl_90 br_90 wl_79 vdd gnd cell_6t
Xbit_r80_c90 bl_90 br_90 wl_80 vdd gnd cell_6t
Xbit_r81_c90 bl_90 br_90 wl_81 vdd gnd cell_6t
Xbit_r82_c90 bl_90 br_90 wl_82 vdd gnd cell_6t
Xbit_r83_c90 bl_90 br_90 wl_83 vdd gnd cell_6t
Xbit_r84_c90 bl_90 br_90 wl_84 vdd gnd cell_6t
Xbit_r85_c90 bl_90 br_90 wl_85 vdd gnd cell_6t
Xbit_r86_c90 bl_90 br_90 wl_86 vdd gnd cell_6t
Xbit_r87_c90 bl_90 br_90 wl_87 vdd gnd cell_6t
Xbit_r88_c90 bl_90 br_90 wl_88 vdd gnd cell_6t
Xbit_r89_c90 bl_90 br_90 wl_89 vdd gnd cell_6t
Xbit_r90_c90 bl_90 br_90 wl_90 vdd gnd cell_6t
Xbit_r91_c90 bl_90 br_90 wl_91 vdd gnd cell_6t
Xbit_r92_c90 bl_90 br_90 wl_92 vdd gnd cell_6t
Xbit_r93_c90 bl_90 br_90 wl_93 vdd gnd cell_6t
Xbit_r94_c90 bl_90 br_90 wl_94 vdd gnd cell_6t
Xbit_r95_c90 bl_90 br_90 wl_95 vdd gnd cell_6t
Xbit_r96_c90 bl_90 br_90 wl_96 vdd gnd cell_6t
Xbit_r97_c90 bl_90 br_90 wl_97 vdd gnd cell_6t
Xbit_r98_c90 bl_90 br_90 wl_98 vdd gnd cell_6t
Xbit_r99_c90 bl_90 br_90 wl_99 vdd gnd cell_6t
Xbit_r100_c90 bl_90 br_90 wl_100 vdd gnd cell_6t
Xbit_r101_c90 bl_90 br_90 wl_101 vdd gnd cell_6t
Xbit_r102_c90 bl_90 br_90 wl_102 vdd gnd cell_6t
Xbit_r103_c90 bl_90 br_90 wl_103 vdd gnd cell_6t
Xbit_r104_c90 bl_90 br_90 wl_104 vdd gnd cell_6t
Xbit_r105_c90 bl_90 br_90 wl_105 vdd gnd cell_6t
Xbit_r106_c90 bl_90 br_90 wl_106 vdd gnd cell_6t
Xbit_r107_c90 bl_90 br_90 wl_107 vdd gnd cell_6t
Xbit_r108_c90 bl_90 br_90 wl_108 vdd gnd cell_6t
Xbit_r109_c90 bl_90 br_90 wl_109 vdd gnd cell_6t
Xbit_r110_c90 bl_90 br_90 wl_110 vdd gnd cell_6t
Xbit_r111_c90 bl_90 br_90 wl_111 vdd gnd cell_6t
Xbit_r112_c90 bl_90 br_90 wl_112 vdd gnd cell_6t
Xbit_r113_c90 bl_90 br_90 wl_113 vdd gnd cell_6t
Xbit_r114_c90 bl_90 br_90 wl_114 vdd gnd cell_6t
Xbit_r115_c90 bl_90 br_90 wl_115 vdd gnd cell_6t
Xbit_r116_c90 bl_90 br_90 wl_116 vdd gnd cell_6t
Xbit_r117_c90 bl_90 br_90 wl_117 vdd gnd cell_6t
Xbit_r118_c90 bl_90 br_90 wl_118 vdd gnd cell_6t
Xbit_r119_c90 bl_90 br_90 wl_119 vdd gnd cell_6t
Xbit_r120_c90 bl_90 br_90 wl_120 vdd gnd cell_6t
Xbit_r121_c90 bl_90 br_90 wl_121 vdd gnd cell_6t
Xbit_r122_c90 bl_90 br_90 wl_122 vdd gnd cell_6t
Xbit_r123_c90 bl_90 br_90 wl_123 vdd gnd cell_6t
Xbit_r124_c90 bl_90 br_90 wl_124 vdd gnd cell_6t
Xbit_r125_c90 bl_90 br_90 wl_125 vdd gnd cell_6t
Xbit_r126_c90 bl_90 br_90 wl_126 vdd gnd cell_6t
Xbit_r127_c90 bl_90 br_90 wl_127 vdd gnd cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd cell_6t
Xbit_r1_c91 bl_91 br_91 wl_1 vdd gnd cell_6t
Xbit_r2_c91 bl_91 br_91 wl_2 vdd gnd cell_6t
Xbit_r3_c91 bl_91 br_91 wl_3 vdd gnd cell_6t
Xbit_r4_c91 bl_91 br_91 wl_4 vdd gnd cell_6t
Xbit_r5_c91 bl_91 br_91 wl_5 vdd gnd cell_6t
Xbit_r6_c91 bl_91 br_91 wl_6 vdd gnd cell_6t
Xbit_r7_c91 bl_91 br_91 wl_7 vdd gnd cell_6t
Xbit_r8_c91 bl_91 br_91 wl_8 vdd gnd cell_6t
Xbit_r9_c91 bl_91 br_91 wl_9 vdd gnd cell_6t
Xbit_r10_c91 bl_91 br_91 wl_10 vdd gnd cell_6t
Xbit_r11_c91 bl_91 br_91 wl_11 vdd gnd cell_6t
Xbit_r12_c91 bl_91 br_91 wl_12 vdd gnd cell_6t
Xbit_r13_c91 bl_91 br_91 wl_13 vdd gnd cell_6t
Xbit_r14_c91 bl_91 br_91 wl_14 vdd gnd cell_6t
Xbit_r15_c91 bl_91 br_91 wl_15 vdd gnd cell_6t
Xbit_r16_c91 bl_91 br_91 wl_16 vdd gnd cell_6t
Xbit_r17_c91 bl_91 br_91 wl_17 vdd gnd cell_6t
Xbit_r18_c91 bl_91 br_91 wl_18 vdd gnd cell_6t
Xbit_r19_c91 bl_91 br_91 wl_19 vdd gnd cell_6t
Xbit_r20_c91 bl_91 br_91 wl_20 vdd gnd cell_6t
Xbit_r21_c91 bl_91 br_91 wl_21 vdd gnd cell_6t
Xbit_r22_c91 bl_91 br_91 wl_22 vdd gnd cell_6t
Xbit_r23_c91 bl_91 br_91 wl_23 vdd gnd cell_6t
Xbit_r24_c91 bl_91 br_91 wl_24 vdd gnd cell_6t
Xbit_r25_c91 bl_91 br_91 wl_25 vdd gnd cell_6t
Xbit_r26_c91 bl_91 br_91 wl_26 vdd gnd cell_6t
Xbit_r27_c91 bl_91 br_91 wl_27 vdd gnd cell_6t
Xbit_r28_c91 bl_91 br_91 wl_28 vdd gnd cell_6t
Xbit_r29_c91 bl_91 br_91 wl_29 vdd gnd cell_6t
Xbit_r30_c91 bl_91 br_91 wl_30 vdd gnd cell_6t
Xbit_r31_c91 bl_91 br_91 wl_31 vdd gnd cell_6t
Xbit_r32_c91 bl_91 br_91 wl_32 vdd gnd cell_6t
Xbit_r33_c91 bl_91 br_91 wl_33 vdd gnd cell_6t
Xbit_r34_c91 bl_91 br_91 wl_34 vdd gnd cell_6t
Xbit_r35_c91 bl_91 br_91 wl_35 vdd gnd cell_6t
Xbit_r36_c91 bl_91 br_91 wl_36 vdd gnd cell_6t
Xbit_r37_c91 bl_91 br_91 wl_37 vdd gnd cell_6t
Xbit_r38_c91 bl_91 br_91 wl_38 vdd gnd cell_6t
Xbit_r39_c91 bl_91 br_91 wl_39 vdd gnd cell_6t
Xbit_r40_c91 bl_91 br_91 wl_40 vdd gnd cell_6t
Xbit_r41_c91 bl_91 br_91 wl_41 vdd gnd cell_6t
Xbit_r42_c91 bl_91 br_91 wl_42 vdd gnd cell_6t
Xbit_r43_c91 bl_91 br_91 wl_43 vdd gnd cell_6t
Xbit_r44_c91 bl_91 br_91 wl_44 vdd gnd cell_6t
Xbit_r45_c91 bl_91 br_91 wl_45 vdd gnd cell_6t
Xbit_r46_c91 bl_91 br_91 wl_46 vdd gnd cell_6t
Xbit_r47_c91 bl_91 br_91 wl_47 vdd gnd cell_6t
Xbit_r48_c91 bl_91 br_91 wl_48 vdd gnd cell_6t
Xbit_r49_c91 bl_91 br_91 wl_49 vdd gnd cell_6t
Xbit_r50_c91 bl_91 br_91 wl_50 vdd gnd cell_6t
Xbit_r51_c91 bl_91 br_91 wl_51 vdd gnd cell_6t
Xbit_r52_c91 bl_91 br_91 wl_52 vdd gnd cell_6t
Xbit_r53_c91 bl_91 br_91 wl_53 vdd gnd cell_6t
Xbit_r54_c91 bl_91 br_91 wl_54 vdd gnd cell_6t
Xbit_r55_c91 bl_91 br_91 wl_55 vdd gnd cell_6t
Xbit_r56_c91 bl_91 br_91 wl_56 vdd gnd cell_6t
Xbit_r57_c91 bl_91 br_91 wl_57 vdd gnd cell_6t
Xbit_r58_c91 bl_91 br_91 wl_58 vdd gnd cell_6t
Xbit_r59_c91 bl_91 br_91 wl_59 vdd gnd cell_6t
Xbit_r60_c91 bl_91 br_91 wl_60 vdd gnd cell_6t
Xbit_r61_c91 bl_91 br_91 wl_61 vdd gnd cell_6t
Xbit_r62_c91 bl_91 br_91 wl_62 vdd gnd cell_6t
Xbit_r63_c91 bl_91 br_91 wl_63 vdd gnd cell_6t
Xbit_r64_c91 bl_91 br_91 wl_64 vdd gnd cell_6t
Xbit_r65_c91 bl_91 br_91 wl_65 vdd gnd cell_6t
Xbit_r66_c91 bl_91 br_91 wl_66 vdd gnd cell_6t
Xbit_r67_c91 bl_91 br_91 wl_67 vdd gnd cell_6t
Xbit_r68_c91 bl_91 br_91 wl_68 vdd gnd cell_6t
Xbit_r69_c91 bl_91 br_91 wl_69 vdd gnd cell_6t
Xbit_r70_c91 bl_91 br_91 wl_70 vdd gnd cell_6t
Xbit_r71_c91 bl_91 br_91 wl_71 vdd gnd cell_6t
Xbit_r72_c91 bl_91 br_91 wl_72 vdd gnd cell_6t
Xbit_r73_c91 bl_91 br_91 wl_73 vdd gnd cell_6t
Xbit_r74_c91 bl_91 br_91 wl_74 vdd gnd cell_6t
Xbit_r75_c91 bl_91 br_91 wl_75 vdd gnd cell_6t
Xbit_r76_c91 bl_91 br_91 wl_76 vdd gnd cell_6t
Xbit_r77_c91 bl_91 br_91 wl_77 vdd gnd cell_6t
Xbit_r78_c91 bl_91 br_91 wl_78 vdd gnd cell_6t
Xbit_r79_c91 bl_91 br_91 wl_79 vdd gnd cell_6t
Xbit_r80_c91 bl_91 br_91 wl_80 vdd gnd cell_6t
Xbit_r81_c91 bl_91 br_91 wl_81 vdd gnd cell_6t
Xbit_r82_c91 bl_91 br_91 wl_82 vdd gnd cell_6t
Xbit_r83_c91 bl_91 br_91 wl_83 vdd gnd cell_6t
Xbit_r84_c91 bl_91 br_91 wl_84 vdd gnd cell_6t
Xbit_r85_c91 bl_91 br_91 wl_85 vdd gnd cell_6t
Xbit_r86_c91 bl_91 br_91 wl_86 vdd gnd cell_6t
Xbit_r87_c91 bl_91 br_91 wl_87 vdd gnd cell_6t
Xbit_r88_c91 bl_91 br_91 wl_88 vdd gnd cell_6t
Xbit_r89_c91 bl_91 br_91 wl_89 vdd gnd cell_6t
Xbit_r90_c91 bl_91 br_91 wl_90 vdd gnd cell_6t
Xbit_r91_c91 bl_91 br_91 wl_91 vdd gnd cell_6t
Xbit_r92_c91 bl_91 br_91 wl_92 vdd gnd cell_6t
Xbit_r93_c91 bl_91 br_91 wl_93 vdd gnd cell_6t
Xbit_r94_c91 bl_91 br_91 wl_94 vdd gnd cell_6t
Xbit_r95_c91 bl_91 br_91 wl_95 vdd gnd cell_6t
Xbit_r96_c91 bl_91 br_91 wl_96 vdd gnd cell_6t
Xbit_r97_c91 bl_91 br_91 wl_97 vdd gnd cell_6t
Xbit_r98_c91 bl_91 br_91 wl_98 vdd gnd cell_6t
Xbit_r99_c91 bl_91 br_91 wl_99 vdd gnd cell_6t
Xbit_r100_c91 bl_91 br_91 wl_100 vdd gnd cell_6t
Xbit_r101_c91 bl_91 br_91 wl_101 vdd gnd cell_6t
Xbit_r102_c91 bl_91 br_91 wl_102 vdd gnd cell_6t
Xbit_r103_c91 bl_91 br_91 wl_103 vdd gnd cell_6t
Xbit_r104_c91 bl_91 br_91 wl_104 vdd gnd cell_6t
Xbit_r105_c91 bl_91 br_91 wl_105 vdd gnd cell_6t
Xbit_r106_c91 bl_91 br_91 wl_106 vdd gnd cell_6t
Xbit_r107_c91 bl_91 br_91 wl_107 vdd gnd cell_6t
Xbit_r108_c91 bl_91 br_91 wl_108 vdd gnd cell_6t
Xbit_r109_c91 bl_91 br_91 wl_109 vdd gnd cell_6t
Xbit_r110_c91 bl_91 br_91 wl_110 vdd gnd cell_6t
Xbit_r111_c91 bl_91 br_91 wl_111 vdd gnd cell_6t
Xbit_r112_c91 bl_91 br_91 wl_112 vdd gnd cell_6t
Xbit_r113_c91 bl_91 br_91 wl_113 vdd gnd cell_6t
Xbit_r114_c91 bl_91 br_91 wl_114 vdd gnd cell_6t
Xbit_r115_c91 bl_91 br_91 wl_115 vdd gnd cell_6t
Xbit_r116_c91 bl_91 br_91 wl_116 vdd gnd cell_6t
Xbit_r117_c91 bl_91 br_91 wl_117 vdd gnd cell_6t
Xbit_r118_c91 bl_91 br_91 wl_118 vdd gnd cell_6t
Xbit_r119_c91 bl_91 br_91 wl_119 vdd gnd cell_6t
Xbit_r120_c91 bl_91 br_91 wl_120 vdd gnd cell_6t
Xbit_r121_c91 bl_91 br_91 wl_121 vdd gnd cell_6t
Xbit_r122_c91 bl_91 br_91 wl_122 vdd gnd cell_6t
Xbit_r123_c91 bl_91 br_91 wl_123 vdd gnd cell_6t
Xbit_r124_c91 bl_91 br_91 wl_124 vdd gnd cell_6t
Xbit_r125_c91 bl_91 br_91 wl_125 vdd gnd cell_6t
Xbit_r126_c91 bl_91 br_91 wl_126 vdd gnd cell_6t
Xbit_r127_c91 bl_91 br_91 wl_127 vdd gnd cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd cell_6t
Xbit_r1_c92 bl_92 br_92 wl_1 vdd gnd cell_6t
Xbit_r2_c92 bl_92 br_92 wl_2 vdd gnd cell_6t
Xbit_r3_c92 bl_92 br_92 wl_3 vdd gnd cell_6t
Xbit_r4_c92 bl_92 br_92 wl_4 vdd gnd cell_6t
Xbit_r5_c92 bl_92 br_92 wl_5 vdd gnd cell_6t
Xbit_r6_c92 bl_92 br_92 wl_6 vdd gnd cell_6t
Xbit_r7_c92 bl_92 br_92 wl_7 vdd gnd cell_6t
Xbit_r8_c92 bl_92 br_92 wl_8 vdd gnd cell_6t
Xbit_r9_c92 bl_92 br_92 wl_9 vdd gnd cell_6t
Xbit_r10_c92 bl_92 br_92 wl_10 vdd gnd cell_6t
Xbit_r11_c92 bl_92 br_92 wl_11 vdd gnd cell_6t
Xbit_r12_c92 bl_92 br_92 wl_12 vdd gnd cell_6t
Xbit_r13_c92 bl_92 br_92 wl_13 vdd gnd cell_6t
Xbit_r14_c92 bl_92 br_92 wl_14 vdd gnd cell_6t
Xbit_r15_c92 bl_92 br_92 wl_15 vdd gnd cell_6t
Xbit_r16_c92 bl_92 br_92 wl_16 vdd gnd cell_6t
Xbit_r17_c92 bl_92 br_92 wl_17 vdd gnd cell_6t
Xbit_r18_c92 bl_92 br_92 wl_18 vdd gnd cell_6t
Xbit_r19_c92 bl_92 br_92 wl_19 vdd gnd cell_6t
Xbit_r20_c92 bl_92 br_92 wl_20 vdd gnd cell_6t
Xbit_r21_c92 bl_92 br_92 wl_21 vdd gnd cell_6t
Xbit_r22_c92 bl_92 br_92 wl_22 vdd gnd cell_6t
Xbit_r23_c92 bl_92 br_92 wl_23 vdd gnd cell_6t
Xbit_r24_c92 bl_92 br_92 wl_24 vdd gnd cell_6t
Xbit_r25_c92 bl_92 br_92 wl_25 vdd gnd cell_6t
Xbit_r26_c92 bl_92 br_92 wl_26 vdd gnd cell_6t
Xbit_r27_c92 bl_92 br_92 wl_27 vdd gnd cell_6t
Xbit_r28_c92 bl_92 br_92 wl_28 vdd gnd cell_6t
Xbit_r29_c92 bl_92 br_92 wl_29 vdd gnd cell_6t
Xbit_r30_c92 bl_92 br_92 wl_30 vdd gnd cell_6t
Xbit_r31_c92 bl_92 br_92 wl_31 vdd gnd cell_6t
Xbit_r32_c92 bl_92 br_92 wl_32 vdd gnd cell_6t
Xbit_r33_c92 bl_92 br_92 wl_33 vdd gnd cell_6t
Xbit_r34_c92 bl_92 br_92 wl_34 vdd gnd cell_6t
Xbit_r35_c92 bl_92 br_92 wl_35 vdd gnd cell_6t
Xbit_r36_c92 bl_92 br_92 wl_36 vdd gnd cell_6t
Xbit_r37_c92 bl_92 br_92 wl_37 vdd gnd cell_6t
Xbit_r38_c92 bl_92 br_92 wl_38 vdd gnd cell_6t
Xbit_r39_c92 bl_92 br_92 wl_39 vdd gnd cell_6t
Xbit_r40_c92 bl_92 br_92 wl_40 vdd gnd cell_6t
Xbit_r41_c92 bl_92 br_92 wl_41 vdd gnd cell_6t
Xbit_r42_c92 bl_92 br_92 wl_42 vdd gnd cell_6t
Xbit_r43_c92 bl_92 br_92 wl_43 vdd gnd cell_6t
Xbit_r44_c92 bl_92 br_92 wl_44 vdd gnd cell_6t
Xbit_r45_c92 bl_92 br_92 wl_45 vdd gnd cell_6t
Xbit_r46_c92 bl_92 br_92 wl_46 vdd gnd cell_6t
Xbit_r47_c92 bl_92 br_92 wl_47 vdd gnd cell_6t
Xbit_r48_c92 bl_92 br_92 wl_48 vdd gnd cell_6t
Xbit_r49_c92 bl_92 br_92 wl_49 vdd gnd cell_6t
Xbit_r50_c92 bl_92 br_92 wl_50 vdd gnd cell_6t
Xbit_r51_c92 bl_92 br_92 wl_51 vdd gnd cell_6t
Xbit_r52_c92 bl_92 br_92 wl_52 vdd gnd cell_6t
Xbit_r53_c92 bl_92 br_92 wl_53 vdd gnd cell_6t
Xbit_r54_c92 bl_92 br_92 wl_54 vdd gnd cell_6t
Xbit_r55_c92 bl_92 br_92 wl_55 vdd gnd cell_6t
Xbit_r56_c92 bl_92 br_92 wl_56 vdd gnd cell_6t
Xbit_r57_c92 bl_92 br_92 wl_57 vdd gnd cell_6t
Xbit_r58_c92 bl_92 br_92 wl_58 vdd gnd cell_6t
Xbit_r59_c92 bl_92 br_92 wl_59 vdd gnd cell_6t
Xbit_r60_c92 bl_92 br_92 wl_60 vdd gnd cell_6t
Xbit_r61_c92 bl_92 br_92 wl_61 vdd gnd cell_6t
Xbit_r62_c92 bl_92 br_92 wl_62 vdd gnd cell_6t
Xbit_r63_c92 bl_92 br_92 wl_63 vdd gnd cell_6t
Xbit_r64_c92 bl_92 br_92 wl_64 vdd gnd cell_6t
Xbit_r65_c92 bl_92 br_92 wl_65 vdd gnd cell_6t
Xbit_r66_c92 bl_92 br_92 wl_66 vdd gnd cell_6t
Xbit_r67_c92 bl_92 br_92 wl_67 vdd gnd cell_6t
Xbit_r68_c92 bl_92 br_92 wl_68 vdd gnd cell_6t
Xbit_r69_c92 bl_92 br_92 wl_69 vdd gnd cell_6t
Xbit_r70_c92 bl_92 br_92 wl_70 vdd gnd cell_6t
Xbit_r71_c92 bl_92 br_92 wl_71 vdd gnd cell_6t
Xbit_r72_c92 bl_92 br_92 wl_72 vdd gnd cell_6t
Xbit_r73_c92 bl_92 br_92 wl_73 vdd gnd cell_6t
Xbit_r74_c92 bl_92 br_92 wl_74 vdd gnd cell_6t
Xbit_r75_c92 bl_92 br_92 wl_75 vdd gnd cell_6t
Xbit_r76_c92 bl_92 br_92 wl_76 vdd gnd cell_6t
Xbit_r77_c92 bl_92 br_92 wl_77 vdd gnd cell_6t
Xbit_r78_c92 bl_92 br_92 wl_78 vdd gnd cell_6t
Xbit_r79_c92 bl_92 br_92 wl_79 vdd gnd cell_6t
Xbit_r80_c92 bl_92 br_92 wl_80 vdd gnd cell_6t
Xbit_r81_c92 bl_92 br_92 wl_81 vdd gnd cell_6t
Xbit_r82_c92 bl_92 br_92 wl_82 vdd gnd cell_6t
Xbit_r83_c92 bl_92 br_92 wl_83 vdd gnd cell_6t
Xbit_r84_c92 bl_92 br_92 wl_84 vdd gnd cell_6t
Xbit_r85_c92 bl_92 br_92 wl_85 vdd gnd cell_6t
Xbit_r86_c92 bl_92 br_92 wl_86 vdd gnd cell_6t
Xbit_r87_c92 bl_92 br_92 wl_87 vdd gnd cell_6t
Xbit_r88_c92 bl_92 br_92 wl_88 vdd gnd cell_6t
Xbit_r89_c92 bl_92 br_92 wl_89 vdd gnd cell_6t
Xbit_r90_c92 bl_92 br_92 wl_90 vdd gnd cell_6t
Xbit_r91_c92 bl_92 br_92 wl_91 vdd gnd cell_6t
Xbit_r92_c92 bl_92 br_92 wl_92 vdd gnd cell_6t
Xbit_r93_c92 bl_92 br_92 wl_93 vdd gnd cell_6t
Xbit_r94_c92 bl_92 br_92 wl_94 vdd gnd cell_6t
Xbit_r95_c92 bl_92 br_92 wl_95 vdd gnd cell_6t
Xbit_r96_c92 bl_92 br_92 wl_96 vdd gnd cell_6t
Xbit_r97_c92 bl_92 br_92 wl_97 vdd gnd cell_6t
Xbit_r98_c92 bl_92 br_92 wl_98 vdd gnd cell_6t
Xbit_r99_c92 bl_92 br_92 wl_99 vdd gnd cell_6t
Xbit_r100_c92 bl_92 br_92 wl_100 vdd gnd cell_6t
Xbit_r101_c92 bl_92 br_92 wl_101 vdd gnd cell_6t
Xbit_r102_c92 bl_92 br_92 wl_102 vdd gnd cell_6t
Xbit_r103_c92 bl_92 br_92 wl_103 vdd gnd cell_6t
Xbit_r104_c92 bl_92 br_92 wl_104 vdd gnd cell_6t
Xbit_r105_c92 bl_92 br_92 wl_105 vdd gnd cell_6t
Xbit_r106_c92 bl_92 br_92 wl_106 vdd gnd cell_6t
Xbit_r107_c92 bl_92 br_92 wl_107 vdd gnd cell_6t
Xbit_r108_c92 bl_92 br_92 wl_108 vdd gnd cell_6t
Xbit_r109_c92 bl_92 br_92 wl_109 vdd gnd cell_6t
Xbit_r110_c92 bl_92 br_92 wl_110 vdd gnd cell_6t
Xbit_r111_c92 bl_92 br_92 wl_111 vdd gnd cell_6t
Xbit_r112_c92 bl_92 br_92 wl_112 vdd gnd cell_6t
Xbit_r113_c92 bl_92 br_92 wl_113 vdd gnd cell_6t
Xbit_r114_c92 bl_92 br_92 wl_114 vdd gnd cell_6t
Xbit_r115_c92 bl_92 br_92 wl_115 vdd gnd cell_6t
Xbit_r116_c92 bl_92 br_92 wl_116 vdd gnd cell_6t
Xbit_r117_c92 bl_92 br_92 wl_117 vdd gnd cell_6t
Xbit_r118_c92 bl_92 br_92 wl_118 vdd gnd cell_6t
Xbit_r119_c92 bl_92 br_92 wl_119 vdd gnd cell_6t
Xbit_r120_c92 bl_92 br_92 wl_120 vdd gnd cell_6t
Xbit_r121_c92 bl_92 br_92 wl_121 vdd gnd cell_6t
Xbit_r122_c92 bl_92 br_92 wl_122 vdd gnd cell_6t
Xbit_r123_c92 bl_92 br_92 wl_123 vdd gnd cell_6t
Xbit_r124_c92 bl_92 br_92 wl_124 vdd gnd cell_6t
Xbit_r125_c92 bl_92 br_92 wl_125 vdd gnd cell_6t
Xbit_r126_c92 bl_92 br_92 wl_126 vdd gnd cell_6t
Xbit_r127_c92 bl_92 br_92 wl_127 vdd gnd cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd cell_6t
Xbit_r1_c93 bl_93 br_93 wl_1 vdd gnd cell_6t
Xbit_r2_c93 bl_93 br_93 wl_2 vdd gnd cell_6t
Xbit_r3_c93 bl_93 br_93 wl_3 vdd gnd cell_6t
Xbit_r4_c93 bl_93 br_93 wl_4 vdd gnd cell_6t
Xbit_r5_c93 bl_93 br_93 wl_5 vdd gnd cell_6t
Xbit_r6_c93 bl_93 br_93 wl_6 vdd gnd cell_6t
Xbit_r7_c93 bl_93 br_93 wl_7 vdd gnd cell_6t
Xbit_r8_c93 bl_93 br_93 wl_8 vdd gnd cell_6t
Xbit_r9_c93 bl_93 br_93 wl_9 vdd gnd cell_6t
Xbit_r10_c93 bl_93 br_93 wl_10 vdd gnd cell_6t
Xbit_r11_c93 bl_93 br_93 wl_11 vdd gnd cell_6t
Xbit_r12_c93 bl_93 br_93 wl_12 vdd gnd cell_6t
Xbit_r13_c93 bl_93 br_93 wl_13 vdd gnd cell_6t
Xbit_r14_c93 bl_93 br_93 wl_14 vdd gnd cell_6t
Xbit_r15_c93 bl_93 br_93 wl_15 vdd gnd cell_6t
Xbit_r16_c93 bl_93 br_93 wl_16 vdd gnd cell_6t
Xbit_r17_c93 bl_93 br_93 wl_17 vdd gnd cell_6t
Xbit_r18_c93 bl_93 br_93 wl_18 vdd gnd cell_6t
Xbit_r19_c93 bl_93 br_93 wl_19 vdd gnd cell_6t
Xbit_r20_c93 bl_93 br_93 wl_20 vdd gnd cell_6t
Xbit_r21_c93 bl_93 br_93 wl_21 vdd gnd cell_6t
Xbit_r22_c93 bl_93 br_93 wl_22 vdd gnd cell_6t
Xbit_r23_c93 bl_93 br_93 wl_23 vdd gnd cell_6t
Xbit_r24_c93 bl_93 br_93 wl_24 vdd gnd cell_6t
Xbit_r25_c93 bl_93 br_93 wl_25 vdd gnd cell_6t
Xbit_r26_c93 bl_93 br_93 wl_26 vdd gnd cell_6t
Xbit_r27_c93 bl_93 br_93 wl_27 vdd gnd cell_6t
Xbit_r28_c93 bl_93 br_93 wl_28 vdd gnd cell_6t
Xbit_r29_c93 bl_93 br_93 wl_29 vdd gnd cell_6t
Xbit_r30_c93 bl_93 br_93 wl_30 vdd gnd cell_6t
Xbit_r31_c93 bl_93 br_93 wl_31 vdd gnd cell_6t
Xbit_r32_c93 bl_93 br_93 wl_32 vdd gnd cell_6t
Xbit_r33_c93 bl_93 br_93 wl_33 vdd gnd cell_6t
Xbit_r34_c93 bl_93 br_93 wl_34 vdd gnd cell_6t
Xbit_r35_c93 bl_93 br_93 wl_35 vdd gnd cell_6t
Xbit_r36_c93 bl_93 br_93 wl_36 vdd gnd cell_6t
Xbit_r37_c93 bl_93 br_93 wl_37 vdd gnd cell_6t
Xbit_r38_c93 bl_93 br_93 wl_38 vdd gnd cell_6t
Xbit_r39_c93 bl_93 br_93 wl_39 vdd gnd cell_6t
Xbit_r40_c93 bl_93 br_93 wl_40 vdd gnd cell_6t
Xbit_r41_c93 bl_93 br_93 wl_41 vdd gnd cell_6t
Xbit_r42_c93 bl_93 br_93 wl_42 vdd gnd cell_6t
Xbit_r43_c93 bl_93 br_93 wl_43 vdd gnd cell_6t
Xbit_r44_c93 bl_93 br_93 wl_44 vdd gnd cell_6t
Xbit_r45_c93 bl_93 br_93 wl_45 vdd gnd cell_6t
Xbit_r46_c93 bl_93 br_93 wl_46 vdd gnd cell_6t
Xbit_r47_c93 bl_93 br_93 wl_47 vdd gnd cell_6t
Xbit_r48_c93 bl_93 br_93 wl_48 vdd gnd cell_6t
Xbit_r49_c93 bl_93 br_93 wl_49 vdd gnd cell_6t
Xbit_r50_c93 bl_93 br_93 wl_50 vdd gnd cell_6t
Xbit_r51_c93 bl_93 br_93 wl_51 vdd gnd cell_6t
Xbit_r52_c93 bl_93 br_93 wl_52 vdd gnd cell_6t
Xbit_r53_c93 bl_93 br_93 wl_53 vdd gnd cell_6t
Xbit_r54_c93 bl_93 br_93 wl_54 vdd gnd cell_6t
Xbit_r55_c93 bl_93 br_93 wl_55 vdd gnd cell_6t
Xbit_r56_c93 bl_93 br_93 wl_56 vdd gnd cell_6t
Xbit_r57_c93 bl_93 br_93 wl_57 vdd gnd cell_6t
Xbit_r58_c93 bl_93 br_93 wl_58 vdd gnd cell_6t
Xbit_r59_c93 bl_93 br_93 wl_59 vdd gnd cell_6t
Xbit_r60_c93 bl_93 br_93 wl_60 vdd gnd cell_6t
Xbit_r61_c93 bl_93 br_93 wl_61 vdd gnd cell_6t
Xbit_r62_c93 bl_93 br_93 wl_62 vdd gnd cell_6t
Xbit_r63_c93 bl_93 br_93 wl_63 vdd gnd cell_6t
Xbit_r64_c93 bl_93 br_93 wl_64 vdd gnd cell_6t
Xbit_r65_c93 bl_93 br_93 wl_65 vdd gnd cell_6t
Xbit_r66_c93 bl_93 br_93 wl_66 vdd gnd cell_6t
Xbit_r67_c93 bl_93 br_93 wl_67 vdd gnd cell_6t
Xbit_r68_c93 bl_93 br_93 wl_68 vdd gnd cell_6t
Xbit_r69_c93 bl_93 br_93 wl_69 vdd gnd cell_6t
Xbit_r70_c93 bl_93 br_93 wl_70 vdd gnd cell_6t
Xbit_r71_c93 bl_93 br_93 wl_71 vdd gnd cell_6t
Xbit_r72_c93 bl_93 br_93 wl_72 vdd gnd cell_6t
Xbit_r73_c93 bl_93 br_93 wl_73 vdd gnd cell_6t
Xbit_r74_c93 bl_93 br_93 wl_74 vdd gnd cell_6t
Xbit_r75_c93 bl_93 br_93 wl_75 vdd gnd cell_6t
Xbit_r76_c93 bl_93 br_93 wl_76 vdd gnd cell_6t
Xbit_r77_c93 bl_93 br_93 wl_77 vdd gnd cell_6t
Xbit_r78_c93 bl_93 br_93 wl_78 vdd gnd cell_6t
Xbit_r79_c93 bl_93 br_93 wl_79 vdd gnd cell_6t
Xbit_r80_c93 bl_93 br_93 wl_80 vdd gnd cell_6t
Xbit_r81_c93 bl_93 br_93 wl_81 vdd gnd cell_6t
Xbit_r82_c93 bl_93 br_93 wl_82 vdd gnd cell_6t
Xbit_r83_c93 bl_93 br_93 wl_83 vdd gnd cell_6t
Xbit_r84_c93 bl_93 br_93 wl_84 vdd gnd cell_6t
Xbit_r85_c93 bl_93 br_93 wl_85 vdd gnd cell_6t
Xbit_r86_c93 bl_93 br_93 wl_86 vdd gnd cell_6t
Xbit_r87_c93 bl_93 br_93 wl_87 vdd gnd cell_6t
Xbit_r88_c93 bl_93 br_93 wl_88 vdd gnd cell_6t
Xbit_r89_c93 bl_93 br_93 wl_89 vdd gnd cell_6t
Xbit_r90_c93 bl_93 br_93 wl_90 vdd gnd cell_6t
Xbit_r91_c93 bl_93 br_93 wl_91 vdd gnd cell_6t
Xbit_r92_c93 bl_93 br_93 wl_92 vdd gnd cell_6t
Xbit_r93_c93 bl_93 br_93 wl_93 vdd gnd cell_6t
Xbit_r94_c93 bl_93 br_93 wl_94 vdd gnd cell_6t
Xbit_r95_c93 bl_93 br_93 wl_95 vdd gnd cell_6t
Xbit_r96_c93 bl_93 br_93 wl_96 vdd gnd cell_6t
Xbit_r97_c93 bl_93 br_93 wl_97 vdd gnd cell_6t
Xbit_r98_c93 bl_93 br_93 wl_98 vdd gnd cell_6t
Xbit_r99_c93 bl_93 br_93 wl_99 vdd gnd cell_6t
Xbit_r100_c93 bl_93 br_93 wl_100 vdd gnd cell_6t
Xbit_r101_c93 bl_93 br_93 wl_101 vdd gnd cell_6t
Xbit_r102_c93 bl_93 br_93 wl_102 vdd gnd cell_6t
Xbit_r103_c93 bl_93 br_93 wl_103 vdd gnd cell_6t
Xbit_r104_c93 bl_93 br_93 wl_104 vdd gnd cell_6t
Xbit_r105_c93 bl_93 br_93 wl_105 vdd gnd cell_6t
Xbit_r106_c93 bl_93 br_93 wl_106 vdd gnd cell_6t
Xbit_r107_c93 bl_93 br_93 wl_107 vdd gnd cell_6t
Xbit_r108_c93 bl_93 br_93 wl_108 vdd gnd cell_6t
Xbit_r109_c93 bl_93 br_93 wl_109 vdd gnd cell_6t
Xbit_r110_c93 bl_93 br_93 wl_110 vdd gnd cell_6t
Xbit_r111_c93 bl_93 br_93 wl_111 vdd gnd cell_6t
Xbit_r112_c93 bl_93 br_93 wl_112 vdd gnd cell_6t
Xbit_r113_c93 bl_93 br_93 wl_113 vdd gnd cell_6t
Xbit_r114_c93 bl_93 br_93 wl_114 vdd gnd cell_6t
Xbit_r115_c93 bl_93 br_93 wl_115 vdd gnd cell_6t
Xbit_r116_c93 bl_93 br_93 wl_116 vdd gnd cell_6t
Xbit_r117_c93 bl_93 br_93 wl_117 vdd gnd cell_6t
Xbit_r118_c93 bl_93 br_93 wl_118 vdd gnd cell_6t
Xbit_r119_c93 bl_93 br_93 wl_119 vdd gnd cell_6t
Xbit_r120_c93 bl_93 br_93 wl_120 vdd gnd cell_6t
Xbit_r121_c93 bl_93 br_93 wl_121 vdd gnd cell_6t
Xbit_r122_c93 bl_93 br_93 wl_122 vdd gnd cell_6t
Xbit_r123_c93 bl_93 br_93 wl_123 vdd gnd cell_6t
Xbit_r124_c93 bl_93 br_93 wl_124 vdd gnd cell_6t
Xbit_r125_c93 bl_93 br_93 wl_125 vdd gnd cell_6t
Xbit_r126_c93 bl_93 br_93 wl_126 vdd gnd cell_6t
Xbit_r127_c93 bl_93 br_93 wl_127 vdd gnd cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd cell_6t
Xbit_r1_c94 bl_94 br_94 wl_1 vdd gnd cell_6t
Xbit_r2_c94 bl_94 br_94 wl_2 vdd gnd cell_6t
Xbit_r3_c94 bl_94 br_94 wl_3 vdd gnd cell_6t
Xbit_r4_c94 bl_94 br_94 wl_4 vdd gnd cell_6t
Xbit_r5_c94 bl_94 br_94 wl_5 vdd gnd cell_6t
Xbit_r6_c94 bl_94 br_94 wl_6 vdd gnd cell_6t
Xbit_r7_c94 bl_94 br_94 wl_7 vdd gnd cell_6t
Xbit_r8_c94 bl_94 br_94 wl_8 vdd gnd cell_6t
Xbit_r9_c94 bl_94 br_94 wl_9 vdd gnd cell_6t
Xbit_r10_c94 bl_94 br_94 wl_10 vdd gnd cell_6t
Xbit_r11_c94 bl_94 br_94 wl_11 vdd gnd cell_6t
Xbit_r12_c94 bl_94 br_94 wl_12 vdd gnd cell_6t
Xbit_r13_c94 bl_94 br_94 wl_13 vdd gnd cell_6t
Xbit_r14_c94 bl_94 br_94 wl_14 vdd gnd cell_6t
Xbit_r15_c94 bl_94 br_94 wl_15 vdd gnd cell_6t
Xbit_r16_c94 bl_94 br_94 wl_16 vdd gnd cell_6t
Xbit_r17_c94 bl_94 br_94 wl_17 vdd gnd cell_6t
Xbit_r18_c94 bl_94 br_94 wl_18 vdd gnd cell_6t
Xbit_r19_c94 bl_94 br_94 wl_19 vdd gnd cell_6t
Xbit_r20_c94 bl_94 br_94 wl_20 vdd gnd cell_6t
Xbit_r21_c94 bl_94 br_94 wl_21 vdd gnd cell_6t
Xbit_r22_c94 bl_94 br_94 wl_22 vdd gnd cell_6t
Xbit_r23_c94 bl_94 br_94 wl_23 vdd gnd cell_6t
Xbit_r24_c94 bl_94 br_94 wl_24 vdd gnd cell_6t
Xbit_r25_c94 bl_94 br_94 wl_25 vdd gnd cell_6t
Xbit_r26_c94 bl_94 br_94 wl_26 vdd gnd cell_6t
Xbit_r27_c94 bl_94 br_94 wl_27 vdd gnd cell_6t
Xbit_r28_c94 bl_94 br_94 wl_28 vdd gnd cell_6t
Xbit_r29_c94 bl_94 br_94 wl_29 vdd gnd cell_6t
Xbit_r30_c94 bl_94 br_94 wl_30 vdd gnd cell_6t
Xbit_r31_c94 bl_94 br_94 wl_31 vdd gnd cell_6t
Xbit_r32_c94 bl_94 br_94 wl_32 vdd gnd cell_6t
Xbit_r33_c94 bl_94 br_94 wl_33 vdd gnd cell_6t
Xbit_r34_c94 bl_94 br_94 wl_34 vdd gnd cell_6t
Xbit_r35_c94 bl_94 br_94 wl_35 vdd gnd cell_6t
Xbit_r36_c94 bl_94 br_94 wl_36 vdd gnd cell_6t
Xbit_r37_c94 bl_94 br_94 wl_37 vdd gnd cell_6t
Xbit_r38_c94 bl_94 br_94 wl_38 vdd gnd cell_6t
Xbit_r39_c94 bl_94 br_94 wl_39 vdd gnd cell_6t
Xbit_r40_c94 bl_94 br_94 wl_40 vdd gnd cell_6t
Xbit_r41_c94 bl_94 br_94 wl_41 vdd gnd cell_6t
Xbit_r42_c94 bl_94 br_94 wl_42 vdd gnd cell_6t
Xbit_r43_c94 bl_94 br_94 wl_43 vdd gnd cell_6t
Xbit_r44_c94 bl_94 br_94 wl_44 vdd gnd cell_6t
Xbit_r45_c94 bl_94 br_94 wl_45 vdd gnd cell_6t
Xbit_r46_c94 bl_94 br_94 wl_46 vdd gnd cell_6t
Xbit_r47_c94 bl_94 br_94 wl_47 vdd gnd cell_6t
Xbit_r48_c94 bl_94 br_94 wl_48 vdd gnd cell_6t
Xbit_r49_c94 bl_94 br_94 wl_49 vdd gnd cell_6t
Xbit_r50_c94 bl_94 br_94 wl_50 vdd gnd cell_6t
Xbit_r51_c94 bl_94 br_94 wl_51 vdd gnd cell_6t
Xbit_r52_c94 bl_94 br_94 wl_52 vdd gnd cell_6t
Xbit_r53_c94 bl_94 br_94 wl_53 vdd gnd cell_6t
Xbit_r54_c94 bl_94 br_94 wl_54 vdd gnd cell_6t
Xbit_r55_c94 bl_94 br_94 wl_55 vdd gnd cell_6t
Xbit_r56_c94 bl_94 br_94 wl_56 vdd gnd cell_6t
Xbit_r57_c94 bl_94 br_94 wl_57 vdd gnd cell_6t
Xbit_r58_c94 bl_94 br_94 wl_58 vdd gnd cell_6t
Xbit_r59_c94 bl_94 br_94 wl_59 vdd gnd cell_6t
Xbit_r60_c94 bl_94 br_94 wl_60 vdd gnd cell_6t
Xbit_r61_c94 bl_94 br_94 wl_61 vdd gnd cell_6t
Xbit_r62_c94 bl_94 br_94 wl_62 vdd gnd cell_6t
Xbit_r63_c94 bl_94 br_94 wl_63 vdd gnd cell_6t
Xbit_r64_c94 bl_94 br_94 wl_64 vdd gnd cell_6t
Xbit_r65_c94 bl_94 br_94 wl_65 vdd gnd cell_6t
Xbit_r66_c94 bl_94 br_94 wl_66 vdd gnd cell_6t
Xbit_r67_c94 bl_94 br_94 wl_67 vdd gnd cell_6t
Xbit_r68_c94 bl_94 br_94 wl_68 vdd gnd cell_6t
Xbit_r69_c94 bl_94 br_94 wl_69 vdd gnd cell_6t
Xbit_r70_c94 bl_94 br_94 wl_70 vdd gnd cell_6t
Xbit_r71_c94 bl_94 br_94 wl_71 vdd gnd cell_6t
Xbit_r72_c94 bl_94 br_94 wl_72 vdd gnd cell_6t
Xbit_r73_c94 bl_94 br_94 wl_73 vdd gnd cell_6t
Xbit_r74_c94 bl_94 br_94 wl_74 vdd gnd cell_6t
Xbit_r75_c94 bl_94 br_94 wl_75 vdd gnd cell_6t
Xbit_r76_c94 bl_94 br_94 wl_76 vdd gnd cell_6t
Xbit_r77_c94 bl_94 br_94 wl_77 vdd gnd cell_6t
Xbit_r78_c94 bl_94 br_94 wl_78 vdd gnd cell_6t
Xbit_r79_c94 bl_94 br_94 wl_79 vdd gnd cell_6t
Xbit_r80_c94 bl_94 br_94 wl_80 vdd gnd cell_6t
Xbit_r81_c94 bl_94 br_94 wl_81 vdd gnd cell_6t
Xbit_r82_c94 bl_94 br_94 wl_82 vdd gnd cell_6t
Xbit_r83_c94 bl_94 br_94 wl_83 vdd gnd cell_6t
Xbit_r84_c94 bl_94 br_94 wl_84 vdd gnd cell_6t
Xbit_r85_c94 bl_94 br_94 wl_85 vdd gnd cell_6t
Xbit_r86_c94 bl_94 br_94 wl_86 vdd gnd cell_6t
Xbit_r87_c94 bl_94 br_94 wl_87 vdd gnd cell_6t
Xbit_r88_c94 bl_94 br_94 wl_88 vdd gnd cell_6t
Xbit_r89_c94 bl_94 br_94 wl_89 vdd gnd cell_6t
Xbit_r90_c94 bl_94 br_94 wl_90 vdd gnd cell_6t
Xbit_r91_c94 bl_94 br_94 wl_91 vdd gnd cell_6t
Xbit_r92_c94 bl_94 br_94 wl_92 vdd gnd cell_6t
Xbit_r93_c94 bl_94 br_94 wl_93 vdd gnd cell_6t
Xbit_r94_c94 bl_94 br_94 wl_94 vdd gnd cell_6t
Xbit_r95_c94 bl_94 br_94 wl_95 vdd gnd cell_6t
Xbit_r96_c94 bl_94 br_94 wl_96 vdd gnd cell_6t
Xbit_r97_c94 bl_94 br_94 wl_97 vdd gnd cell_6t
Xbit_r98_c94 bl_94 br_94 wl_98 vdd gnd cell_6t
Xbit_r99_c94 bl_94 br_94 wl_99 vdd gnd cell_6t
Xbit_r100_c94 bl_94 br_94 wl_100 vdd gnd cell_6t
Xbit_r101_c94 bl_94 br_94 wl_101 vdd gnd cell_6t
Xbit_r102_c94 bl_94 br_94 wl_102 vdd gnd cell_6t
Xbit_r103_c94 bl_94 br_94 wl_103 vdd gnd cell_6t
Xbit_r104_c94 bl_94 br_94 wl_104 vdd gnd cell_6t
Xbit_r105_c94 bl_94 br_94 wl_105 vdd gnd cell_6t
Xbit_r106_c94 bl_94 br_94 wl_106 vdd gnd cell_6t
Xbit_r107_c94 bl_94 br_94 wl_107 vdd gnd cell_6t
Xbit_r108_c94 bl_94 br_94 wl_108 vdd gnd cell_6t
Xbit_r109_c94 bl_94 br_94 wl_109 vdd gnd cell_6t
Xbit_r110_c94 bl_94 br_94 wl_110 vdd gnd cell_6t
Xbit_r111_c94 bl_94 br_94 wl_111 vdd gnd cell_6t
Xbit_r112_c94 bl_94 br_94 wl_112 vdd gnd cell_6t
Xbit_r113_c94 bl_94 br_94 wl_113 vdd gnd cell_6t
Xbit_r114_c94 bl_94 br_94 wl_114 vdd gnd cell_6t
Xbit_r115_c94 bl_94 br_94 wl_115 vdd gnd cell_6t
Xbit_r116_c94 bl_94 br_94 wl_116 vdd gnd cell_6t
Xbit_r117_c94 bl_94 br_94 wl_117 vdd gnd cell_6t
Xbit_r118_c94 bl_94 br_94 wl_118 vdd gnd cell_6t
Xbit_r119_c94 bl_94 br_94 wl_119 vdd gnd cell_6t
Xbit_r120_c94 bl_94 br_94 wl_120 vdd gnd cell_6t
Xbit_r121_c94 bl_94 br_94 wl_121 vdd gnd cell_6t
Xbit_r122_c94 bl_94 br_94 wl_122 vdd gnd cell_6t
Xbit_r123_c94 bl_94 br_94 wl_123 vdd gnd cell_6t
Xbit_r124_c94 bl_94 br_94 wl_124 vdd gnd cell_6t
Xbit_r125_c94 bl_94 br_94 wl_125 vdd gnd cell_6t
Xbit_r126_c94 bl_94 br_94 wl_126 vdd gnd cell_6t
Xbit_r127_c94 bl_94 br_94 wl_127 vdd gnd cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd cell_6t
Xbit_r1_c95 bl_95 br_95 wl_1 vdd gnd cell_6t
Xbit_r2_c95 bl_95 br_95 wl_2 vdd gnd cell_6t
Xbit_r3_c95 bl_95 br_95 wl_3 vdd gnd cell_6t
Xbit_r4_c95 bl_95 br_95 wl_4 vdd gnd cell_6t
Xbit_r5_c95 bl_95 br_95 wl_5 vdd gnd cell_6t
Xbit_r6_c95 bl_95 br_95 wl_6 vdd gnd cell_6t
Xbit_r7_c95 bl_95 br_95 wl_7 vdd gnd cell_6t
Xbit_r8_c95 bl_95 br_95 wl_8 vdd gnd cell_6t
Xbit_r9_c95 bl_95 br_95 wl_9 vdd gnd cell_6t
Xbit_r10_c95 bl_95 br_95 wl_10 vdd gnd cell_6t
Xbit_r11_c95 bl_95 br_95 wl_11 vdd gnd cell_6t
Xbit_r12_c95 bl_95 br_95 wl_12 vdd gnd cell_6t
Xbit_r13_c95 bl_95 br_95 wl_13 vdd gnd cell_6t
Xbit_r14_c95 bl_95 br_95 wl_14 vdd gnd cell_6t
Xbit_r15_c95 bl_95 br_95 wl_15 vdd gnd cell_6t
Xbit_r16_c95 bl_95 br_95 wl_16 vdd gnd cell_6t
Xbit_r17_c95 bl_95 br_95 wl_17 vdd gnd cell_6t
Xbit_r18_c95 bl_95 br_95 wl_18 vdd gnd cell_6t
Xbit_r19_c95 bl_95 br_95 wl_19 vdd gnd cell_6t
Xbit_r20_c95 bl_95 br_95 wl_20 vdd gnd cell_6t
Xbit_r21_c95 bl_95 br_95 wl_21 vdd gnd cell_6t
Xbit_r22_c95 bl_95 br_95 wl_22 vdd gnd cell_6t
Xbit_r23_c95 bl_95 br_95 wl_23 vdd gnd cell_6t
Xbit_r24_c95 bl_95 br_95 wl_24 vdd gnd cell_6t
Xbit_r25_c95 bl_95 br_95 wl_25 vdd gnd cell_6t
Xbit_r26_c95 bl_95 br_95 wl_26 vdd gnd cell_6t
Xbit_r27_c95 bl_95 br_95 wl_27 vdd gnd cell_6t
Xbit_r28_c95 bl_95 br_95 wl_28 vdd gnd cell_6t
Xbit_r29_c95 bl_95 br_95 wl_29 vdd gnd cell_6t
Xbit_r30_c95 bl_95 br_95 wl_30 vdd gnd cell_6t
Xbit_r31_c95 bl_95 br_95 wl_31 vdd gnd cell_6t
Xbit_r32_c95 bl_95 br_95 wl_32 vdd gnd cell_6t
Xbit_r33_c95 bl_95 br_95 wl_33 vdd gnd cell_6t
Xbit_r34_c95 bl_95 br_95 wl_34 vdd gnd cell_6t
Xbit_r35_c95 bl_95 br_95 wl_35 vdd gnd cell_6t
Xbit_r36_c95 bl_95 br_95 wl_36 vdd gnd cell_6t
Xbit_r37_c95 bl_95 br_95 wl_37 vdd gnd cell_6t
Xbit_r38_c95 bl_95 br_95 wl_38 vdd gnd cell_6t
Xbit_r39_c95 bl_95 br_95 wl_39 vdd gnd cell_6t
Xbit_r40_c95 bl_95 br_95 wl_40 vdd gnd cell_6t
Xbit_r41_c95 bl_95 br_95 wl_41 vdd gnd cell_6t
Xbit_r42_c95 bl_95 br_95 wl_42 vdd gnd cell_6t
Xbit_r43_c95 bl_95 br_95 wl_43 vdd gnd cell_6t
Xbit_r44_c95 bl_95 br_95 wl_44 vdd gnd cell_6t
Xbit_r45_c95 bl_95 br_95 wl_45 vdd gnd cell_6t
Xbit_r46_c95 bl_95 br_95 wl_46 vdd gnd cell_6t
Xbit_r47_c95 bl_95 br_95 wl_47 vdd gnd cell_6t
Xbit_r48_c95 bl_95 br_95 wl_48 vdd gnd cell_6t
Xbit_r49_c95 bl_95 br_95 wl_49 vdd gnd cell_6t
Xbit_r50_c95 bl_95 br_95 wl_50 vdd gnd cell_6t
Xbit_r51_c95 bl_95 br_95 wl_51 vdd gnd cell_6t
Xbit_r52_c95 bl_95 br_95 wl_52 vdd gnd cell_6t
Xbit_r53_c95 bl_95 br_95 wl_53 vdd gnd cell_6t
Xbit_r54_c95 bl_95 br_95 wl_54 vdd gnd cell_6t
Xbit_r55_c95 bl_95 br_95 wl_55 vdd gnd cell_6t
Xbit_r56_c95 bl_95 br_95 wl_56 vdd gnd cell_6t
Xbit_r57_c95 bl_95 br_95 wl_57 vdd gnd cell_6t
Xbit_r58_c95 bl_95 br_95 wl_58 vdd gnd cell_6t
Xbit_r59_c95 bl_95 br_95 wl_59 vdd gnd cell_6t
Xbit_r60_c95 bl_95 br_95 wl_60 vdd gnd cell_6t
Xbit_r61_c95 bl_95 br_95 wl_61 vdd gnd cell_6t
Xbit_r62_c95 bl_95 br_95 wl_62 vdd gnd cell_6t
Xbit_r63_c95 bl_95 br_95 wl_63 vdd gnd cell_6t
Xbit_r64_c95 bl_95 br_95 wl_64 vdd gnd cell_6t
Xbit_r65_c95 bl_95 br_95 wl_65 vdd gnd cell_6t
Xbit_r66_c95 bl_95 br_95 wl_66 vdd gnd cell_6t
Xbit_r67_c95 bl_95 br_95 wl_67 vdd gnd cell_6t
Xbit_r68_c95 bl_95 br_95 wl_68 vdd gnd cell_6t
Xbit_r69_c95 bl_95 br_95 wl_69 vdd gnd cell_6t
Xbit_r70_c95 bl_95 br_95 wl_70 vdd gnd cell_6t
Xbit_r71_c95 bl_95 br_95 wl_71 vdd gnd cell_6t
Xbit_r72_c95 bl_95 br_95 wl_72 vdd gnd cell_6t
Xbit_r73_c95 bl_95 br_95 wl_73 vdd gnd cell_6t
Xbit_r74_c95 bl_95 br_95 wl_74 vdd gnd cell_6t
Xbit_r75_c95 bl_95 br_95 wl_75 vdd gnd cell_6t
Xbit_r76_c95 bl_95 br_95 wl_76 vdd gnd cell_6t
Xbit_r77_c95 bl_95 br_95 wl_77 vdd gnd cell_6t
Xbit_r78_c95 bl_95 br_95 wl_78 vdd gnd cell_6t
Xbit_r79_c95 bl_95 br_95 wl_79 vdd gnd cell_6t
Xbit_r80_c95 bl_95 br_95 wl_80 vdd gnd cell_6t
Xbit_r81_c95 bl_95 br_95 wl_81 vdd gnd cell_6t
Xbit_r82_c95 bl_95 br_95 wl_82 vdd gnd cell_6t
Xbit_r83_c95 bl_95 br_95 wl_83 vdd gnd cell_6t
Xbit_r84_c95 bl_95 br_95 wl_84 vdd gnd cell_6t
Xbit_r85_c95 bl_95 br_95 wl_85 vdd gnd cell_6t
Xbit_r86_c95 bl_95 br_95 wl_86 vdd gnd cell_6t
Xbit_r87_c95 bl_95 br_95 wl_87 vdd gnd cell_6t
Xbit_r88_c95 bl_95 br_95 wl_88 vdd gnd cell_6t
Xbit_r89_c95 bl_95 br_95 wl_89 vdd gnd cell_6t
Xbit_r90_c95 bl_95 br_95 wl_90 vdd gnd cell_6t
Xbit_r91_c95 bl_95 br_95 wl_91 vdd gnd cell_6t
Xbit_r92_c95 bl_95 br_95 wl_92 vdd gnd cell_6t
Xbit_r93_c95 bl_95 br_95 wl_93 vdd gnd cell_6t
Xbit_r94_c95 bl_95 br_95 wl_94 vdd gnd cell_6t
Xbit_r95_c95 bl_95 br_95 wl_95 vdd gnd cell_6t
Xbit_r96_c95 bl_95 br_95 wl_96 vdd gnd cell_6t
Xbit_r97_c95 bl_95 br_95 wl_97 vdd gnd cell_6t
Xbit_r98_c95 bl_95 br_95 wl_98 vdd gnd cell_6t
Xbit_r99_c95 bl_95 br_95 wl_99 vdd gnd cell_6t
Xbit_r100_c95 bl_95 br_95 wl_100 vdd gnd cell_6t
Xbit_r101_c95 bl_95 br_95 wl_101 vdd gnd cell_6t
Xbit_r102_c95 bl_95 br_95 wl_102 vdd gnd cell_6t
Xbit_r103_c95 bl_95 br_95 wl_103 vdd gnd cell_6t
Xbit_r104_c95 bl_95 br_95 wl_104 vdd gnd cell_6t
Xbit_r105_c95 bl_95 br_95 wl_105 vdd gnd cell_6t
Xbit_r106_c95 bl_95 br_95 wl_106 vdd gnd cell_6t
Xbit_r107_c95 bl_95 br_95 wl_107 vdd gnd cell_6t
Xbit_r108_c95 bl_95 br_95 wl_108 vdd gnd cell_6t
Xbit_r109_c95 bl_95 br_95 wl_109 vdd gnd cell_6t
Xbit_r110_c95 bl_95 br_95 wl_110 vdd gnd cell_6t
Xbit_r111_c95 bl_95 br_95 wl_111 vdd gnd cell_6t
Xbit_r112_c95 bl_95 br_95 wl_112 vdd gnd cell_6t
Xbit_r113_c95 bl_95 br_95 wl_113 vdd gnd cell_6t
Xbit_r114_c95 bl_95 br_95 wl_114 vdd gnd cell_6t
Xbit_r115_c95 bl_95 br_95 wl_115 vdd gnd cell_6t
Xbit_r116_c95 bl_95 br_95 wl_116 vdd gnd cell_6t
Xbit_r117_c95 bl_95 br_95 wl_117 vdd gnd cell_6t
Xbit_r118_c95 bl_95 br_95 wl_118 vdd gnd cell_6t
Xbit_r119_c95 bl_95 br_95 wl_119 vdd gnd cell_6t
Xbit_r120_c95 bl_95 br_95 wl_120 vdd gnd cell_6t
Xbit_r121_c95 bl_95 br_95 wl_121 vdd gnd cell_6t
Xbit_r122_c95 bl_95 br_95 wl_122 vdd gnd cell_6t
Xbit_r123_c95 bl_95 br_95 wl_123 vdd gnd cell_6t
Xbit_r124_c95 bl_95 br_95 wl_124 vdd gnd cell_6t
Xbit_r125_c95 bl_95 br_95 wl_125 vdd gnd cell_6t
Xbit_r126_c95 bl_95 br_95 wl_126 vdd gnd cell_6t
Xbit_r127_c95 bl_95 br_95 wl_127 vdd gnd cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd cell_6t
Xbit_r1_c96 bl_96 br_96 wl_1 vdd gnd cell_6t
Xbit_r2_c96 bl_96 br_96 wl_2 vdd gnd cell_6t
Xbit_r3_c96 bl_96 br_96 wl_3 vdd gnd cell_6t
Xbit_r4_c96 bl_96 br_96 wl_4 vdd gnd cell_6t
Xbit_r5_c96 bl_96 br_96 wl_5 vdd gnd cell_6t
Xbit_r6_c96 bl_96 br_96 wl_6 vdd gnd cell_6t
Xbit_r7_c96 bl_96 br_96 wl_7 vdd gnd cell_6t
Xbit_r8_c96 bl_96 br_96 wl_8 vdd gnd cell_6t
Xbit_r9_c96 bl_96 br_96 wl_9 vdd gnd cell_6t
Xbit_r10_c96 bl_96 br_96 wl_10 vdd gnd cell_6t
Xbit_r11_c96 bl_96 br_96 wl_11 vdd gnd cell_6t
Xbit_r12_c96 bl_96 br_96 wl_12 vdd gnd cell_6t
Xbit_r13_c96 bl_96 br_96 wl_13 vdd gnd cell_6t
Xbit_r14_c96 bl_96 br_96 wl_14 vdd gnd cell_6t
Xbit_r15_c96 bl_96 br_96 wl_15 vdd gnd cell_6t
Xbit_r16_c96 bl_96 br_96 wl_16 vdd gnd cell_6t
Xbit_r17_c96 bl_96 br_96 wl_17 vdd gnd cell_6t
Xbit_r18_c96 bl_96 br_96 wl_18 vdd gnd cell_6t
Xbit_r19_c96 bl_96 br_96 wl_19 vdd gnd cell_6t
Xbit_r20_c96 bl_96 br_96 wl_20 vdd gnd cell_6t
Xbit_r21_c96 bl_96 br_96 wl_21 vdd gnd cell_6t
Xbit_r22_c96 bl_96 br_96 wl_22 vdd gnd cell_6t
Xbit_r23_c96 bl_96 br_96 wl_23 vdd gnd cell_6t
Xbit_r24_c96 bl_96 br_96 wl_24 vdd gnd cell_6t
Xbit_r25_c96 bl_96 br_96 wl_25 vdd gnd cell_6t
Xbit_r26_c96 bl_96 br_96 wl_26 vdd gnd cell_6t
Xbit_r27_c96 bl_96 br_96 wl_27 vdd gnd cell_6t
Xbit_r28_c96 bl_96 br_96 wl_28 vdd gnd cell_6t
Xbit_r29_c96 bl_96 br_96 wl_29 vdd gnd cell_6t
Xbit_r30_c96 bl_96 br_96 wl_30 vdd gnd cell_6t
Xbit_r31_c96 bl_96 br_96 wl_31 vdd gnd cell_6t
Xbit_r32_c96 bl_96 br_96 wl_32 vdd gnd cell_6t
Xbit_r33_c96 bl_96 br_96 wl_33 vdd gnd cell_6t
Xbit_r34_c96 bl_96 br_96 wl_34 vdd gnd cell_6t
Xbit_r35_c96 bl_96 br_96 wl_35 vdd gnd cell_6t
Xbit_r36_c96 bl_96 br_96 wl_36 vdd gnd cell_6t
Xbit_r37_c96 bl_96 br_96 wl_37 vdd gnd cell_6t
Xbit_r38_c96 bl_96 br_96 wl_38 vdd gnd cell_6t
Xbit_r39_c96 bl_96 br_96 wl_39 vdd gnd cell_6t
Xbit_r40_c96 bl_96 br_96 wl_40 vdd gnd cell_6t
Xbit_r41_c96 bl_96 br_96 wl_41 vdd gnd cell_6t
Xbit_r42_c96 bl_96 br_96 wl_42 vdd gnd cell_6t
Xbit_r43_c96 bl_96 br_96 wl_43 vdd gnd cell_6t
Xbit_r44_c96 bl_96 br_96 wl_44 vdd gnd cell_6t
Xbit_r45_c96 bl_96 br_96 wl_45 vdd gnd cell_6t
Xbit_r46_c96 bl_96 br_96 wl_46 vdd gnd cell_6t
Xbit_r47_c96 bl_96 br_96 wl_47 vdd gnd cell_6t
Xbit_r48_c96 bl_96 br_96 wl_48 vdd gnd cell_6t
Xbit_r49_c96 bl_96 br_96 wl_49 vdd gnd cell_6t
Xbit_r50_c96 bl_96 br_96 wl_50 vdd gnd cell_6t
Xbit_r51_c96 bl_96 br_96 wl_51 vdd gnd cell_6t
Xbit_r52_c96 bl_96 br_96 wl_52 vdd gnd cell_6t
Xbit_r53_c96 bl_96 br_96 wl_53 vdd gnd cell_6t
Xbit_r54_c96 bl_96 br_96 wl_54 vdd gnd cell_6t
Xbit_r55_c96 bl_96 br_96 wl_55 vdd gnd cell_6t
Xbit_r56_c96 bl_96 br_96 wl_56 vdd gnd cell_6t
Xbit_r57_c96 bl_96 br_96 wl_57 vdd gnd cell_6t
Xbit_r58_c96 bl_96 br_96 wl_58 vdd gnd cell_6t
Xbit_r59_c96 bl_96 br_96 wl_59 vdd gnd cell_6t
Xbit_r60_c96 bl_96 br_96 wl_60 vdd gnd cell_6t
Xbit_r61_c96 bl_96 br_96 wl_61 vdd gnd cell_6t
Xbit_r62_c96 bl_96 br_96 wl_62 vdd gnd cell_6t
Xbit_r63_c96 bl_96 br_96 wl_63 vdd gnd cell_6t
Xbit_r64_c96 bl_96 br_96 wl_64 vdd gnd cell_6t
Xbit_r65_c96 bl_96 br_96 wl_65 vdd gnd cell_6t
Xbit_r66_c96 bl_96 br_96 wl_66 vdd gnd cell_6t
Xbit_r67_c96 bl_96 br_96 wl_67 vdd gnd cell_6t
Xbit_r68_c96 bl_96 br_96 wl_68 vdd gnd cell_6t
Xbit_r69_c96 bl_96 br_96 wl_69 vdd gnd cell_6t
Xbit_r70_c96 bl_96 br_96 wl_70 vdd gnd cell_6t
Xbit_r71_c96 bl_96 br_96 wl_71 vdd gnd cell_6t
Xbit_r72_c96 bl_96 br_96 wl_72 vdd gnd cell_6t
Xbit_r73_c96 bl_96 br_96 wl_73 vdd gnd cell_6t
Xbit_r74_c96 bl_96 br_96 wl_74 vdd gnd cell_6t
Xbit_r75_c96 bl_96 br_96 wl_75 vdd gnd cell_6t
Xbit_r76_c96 bl_96 br_96 wl_76 vdd gnd cell_6t
Xbit_r77_c96 bl_96 br_96 wl_77 vdd gnd cell_6t
Xbit_r78_c96 bl_96 br_96 wl_78 vdd gnd cell_6t
Xbit_r79_c96 bl_96 br_96 wl_79 vdd gnd cell_6t
Xbit_r80_c96 bl_96 br_96 wl_80 vdd gnd cell_6t
Xbit_r81_c96 bl_96 br_96 wl_81 vdd gnd cell_6t
Xbit_r82_c96 bl_96 br_96 wl_82 vdd gnd cell_6t
Xbit_r83_c96 bl_96 br_96 wl_83 vdd gnd cell_6t
Xbit_r84_c96 bl_96 br_96 wl_84 vdd gnd cell_6t
Xbit_r85_c96 bl_96 br_96 wl_85 vdd gnd cell_6t
Xbit_r86_c96 bl_96 br_96 wl_86 vdd gnd cell_6t
Xbit_r87_c96 bl_96 br_96 wl_87 vdd gnd cell_6t
Xbit_r88_c96 bl_96 br_96 wl_88 vdd gnd cell_6t
Xbit_r89_c96 bl_96 br_96 wl_89 vdd gnd cell_6t
Xbit_r90_c96 bl_96 br_96 wl_90 vdd gnd cell_6t
Xbit_r91_c96 bl_96 br_96 wl_91 vdd gnd cell_6t
Xbit_r92_c96 bl_96 br_96 wl_92 vdd gnd cell_6t
Xbit_r93_c96 bl_96 br_96 wl_93 vdd gnd cell_6t
Xbit_r94_c96 bl_96 br_96 wl_94 vdd gnd cell_6t
Xbit_r95_c96 bl_96 br_96 wl_95 vdd gnd cell_6t
Xbit_r96_c96 bl_96 br_96 wl_96 vdd gnd cell_6t
Xbit_r97_c96 bl_96 br_96 wl_97 vdd gnd cell_6t
Xbit_r98_c96 bl_96 br_96 wl_98 vdd gnd cell_6t
Xbit_r99_c96 bl_96 br_96 wl_99 vdd gnd cell_6t
Xbit_r100_c96 bl_96 br_96 wl_100 vdd gnd cell_6t
Xbit_r101_c96 bl_96 br_96 wl_101 vdd gnd cell_6t
Xbit_r102_c96 bl_96 br_96 wl_102 vdd gnd cell_6t
Xbit_r103_c96 bl_96 br_96 wl_103 vdd gnd cell_6t
Xbit_r104_c96 bl_96 br_96 wl_104 vdd gnd cell_6t
Xbit_r105_c96 bl_96 br_96 wl_105 vdd gnd cell_6t
Xbit_r106_c96 bl_96 br_96 wl_106 vdd gnd cell_6t
Xbit_r107_c96 bl_96 br_96 wl_107 vdd gnd cell_6t
Xbit_r108_c96 bl_96 br_96 wl_108 vdd gnd cell_6t
Xbit_r109_c96 bl_96 br_96 wl_109 vdd gnd cell_6t
Xbit_r110_c96 bl_96 br_96 wl_110 vdd gnd cell_6t
Xbit_r111_c96 bl_96 br_96 wl_111 vdd gnd cell_6t
Xbit_r112_c96 bl_96 br_96 wl_112 vdd gnd cell_6t
Xbit_r113_c96 bl_96 br_96 wl_113 vdd gnd cell_6t
Xbit_r114_c96 bl_96 br_96 wl_114 vdd gnd cell_6t
Xbit_r115_c96 bl_96 br_96 wl_115 vdd gnd cell_6t
Xbit_r116_c96 bl_96 br_96 wl_116 vdd gnd cell_6t
Xbit_r117_c96 bl_96 br_96 wl_117 vdd gnd cell_6t
Xbit_r118_c96 bl_96 br_96 wl_118 vdd gnd cell_6t
Xbit_r119_c96 bl_96 br_96 wl_119 vdd gnd cell_6t
Xbit_r120_c96 bl_96 br_96 wl_120 vdd gnd cell_6t
Xbit_r121_c96 bl_96 br_96 wl_121 vdd gnd cell_6t
Xbit_r122_c96 bl_96 br_96 wl_122 vdd gnd cell_6t
Xbit_r123_c96 bl_96 br_96 wl_123 vdd gnd cell_6t
Xbit_r124_c96 bl_96 br_96 wl_124 vdd gnd cell_6t
Xbit_r125_c96 bl_96 br_96 wl_125 vdd gnd cell_6t
Xbit_r126_c96 bl_96 br_96 wl_126 vdd gnd cell_6t
Xbit_r127_c96 bl_96 br_96 wl_127 vdd gnd cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd cell_6t
Xbit_r1_c97 bl_97 br_97 wl_1 vdd gnd cell_6t
Xbit_r2_c97 bl_97 br_97 wl_2 vdd gnd cell_6t
Xbit_r3_c97 bl_97 br_97 wl_3 vdd gnd cell_6t
Xbit_r4_c97 bl_97 br_97 wl_4 vdd gnd cell_6t
Xbit_r5_c97 bl_97 br_97 wl_5 vdd gnd cell_6t
Xbit_r6_c97 bl_97 br_97 wl_6 vdd gnd cell_6t
Xbit_r7_c97 bl_97 br_97 wl_7 vdd gnd cell_6t
Xbit_r8_c97 bl_97 br_97 wl_8 vdd gnd cell_6t
Xbit_r9_c97 bl_97 br_97 wl_9 vdd gnd cell_6t
Xbit_r10_c97 bl_97 br_97 wl_10 vdd gnd cell_6t
Xbit_r11_c97 bl_97 br_97 wl_11 vdd gnd cell_6t
Xbit_r12_c97 bl_97 br_97 wl_12 vdd gnd cell_6t
Xbit_r13_c97 bl_97 br_97 wl_13 vdd gnd cell_6t
Xbit_r14_c97 bl_97 br_97 wl_14 vdd gnd cell_6t
Xbit_r15_c97 bl_97 br_97 wl_15 vdd gnd cell_6t
Xbit_r16_c97 bl_97 br_97 wl_16 vdd gnd cell_6t
Xbit_r17_c97 bl_97 br_97 wl_17 vdd gnd cell_6t
Xbit_r18_c97 bl_97 br_97 wl_18 vdd gnd cell_6t
Xbit_r19_c97 bl_97 br_97 wl_19 vdd gnd cell_6t
Xbit_r20_c97 bl_97 br_97 wl_20 vdd gnd cell_6t
Xbit_r21_c97 bl_97 br_97 wl_21 vdd gnd cell_6t
Xbit_r22_c97 bl_97 br_97 wl_22 vdd gnd cell_6t
Xbit_r23_c97 bl_97 br_97 wl_23 vdd gnd cell_6t
Xbit_r24_c97 bl_97 br_97 wl_24 vdd gnd cell_6t
Xbit_r25_c97 bl_97 br_97 wl_25 vdd gnd cell_6t
Xbit_r26_c97 bl_97 br_97 wl_26 vdd gnd cell_6t
Xbit_r27_c97 bl_97 br_97 wl_27 vdd gnd cell_6t
Xbit_r28_c97 bl_97 br_97 wl_28 vdd gnd cell_6t
Xbit_r29_c97 bl_97 br_97 wl_29 vdd gnd cell_6t
Xbit_r30_c97 bl_97 br_97 wl_30 vdd gnd cell_6t
Xbit_r31_c97 bl_97 br_97 wl_31 vdd gnd cell_6t
Xbit_r32_c97 bl_97 br_97 wl_32 vdd gnd cell_6t
Xbit_r33_c97 bl_97 br_97 wl_33 vdd gnd cell_6t
Xbit_r34_c97 bl_97 br_97 wl_34 vdd gnd cell_6t
Xbit_r35_c97 bl_97 br_97 wl_35 vdd gnd cell_6t
Xbit_r36_c97 bl_97 br_97 wl_36 vdd gnd cell_6t
Xbit_r37_c97 bl_97 br_97 wl_37 vdd gnd cell_6t
Xbit_r38_c97 bl_97 br_97 wl_38 vdd gnd cell_6t
Xbit_r39_c97 bl_97 br_97 wl_39 vdd gnd cell_6t
Xbit_r40_c97 bl_97 br_97 wl_40 vdd gnd cell_6t
Xbit_r41_c97 bl_97 br_97 wl_41 vdd gnd cell_6t
Xbit_r42_c97 bl_97 br_97 wl_42 vdd gnd cell_6t
Xbit_r43_c97 bl_97 br_97 wl_43 vdd gnd cell_6t
Xbit_r44_c97 bl_97 br_97 wl_44 vdd gnd cell_6t
Xbit_r45_c97 bl_97 br_97 wl_45 vdd gnd cell_6t
Xbit_r46_c97 bl_97 br_97 wl_46 vdd gnd cell_6t
Xbit_r47_c97 bl_97 br_97 wl_47 vdd gnd cell_6t
Xbit_r48_c97 bl_97 br_97 wl_48 vdd gnd cell_6t
Xbit_r49_c97 bl_97 br_97 wl_49 vdd gnd cell_6t
Xbit_r50_c97 bl_97 br_97 wl_50 vdd gnd cell_6t
Xbit_r51_c97 bl_97 br_97 wl_51 vdd gnd cell_6t
Xbit_r52_c97 bl_97 br_97 wl_52 vdd gnd cell_6t
Xbit_r53_c97 bl_97 br_97 wl_53 vdd gnd cell_6t
Xbit_r54_c97 bl_97 br_97 wl_54 vdd gnd cell_6t
Xbit_r55_c97 bl_97 br_97 wl_55 vdd gnd cell_6t
Xbit_r56_c97 bl_97 br_97 wl_56 vdd gnd cell_6t
Xbit_r57_c97 bl_97 br_97 wl_57 vdd gnd cell_6t
Xbit_r58_c97 bl_97 br_97 wl_58 vdd gnd cell_6t
Xbit_r59_c97 bl_97 br_97 wl_59 vdd gnd cell_6t
Xbit_r60_c97 bl_97 br_97 wl_60 vdd gnd cell_6t
Xbit_r61_c97 bl_97 br_97 wl_61 vdd gnd cell_6t
Xbit_r62_c97 bl_97 br_97 wl_62 vdd gnd cell_6t
Xbit_r63_c97 bl_97 br_97 wl_63 vdd gnd cell_6t
Xbit_r64_c97 bl_97 br_97 wl_64 vdd gnd cell_6t
Xbit_r65_c97 bl_97 br_97 wl_65 vdd gnd cell_6t
Xbit_r66_c97 bl_97 br_97 wl_66 vdd gnd cell_6t
Xbit_r67_c97 bl_97 br_97 wl_67 vdd gnd cell_6t
Xbit_r68_c97 bl_97 br_97 wl_68 vdd gnd cell_6t
Xbit_r69_c97 bl_97 br_97 wl_69 vdd gnd cell_6t
Xbit_r70_c97 bl_97 br_97 wl_70 vdd gnd cell_6t
Xbit_r71_c97 bl_97 br_97 wl_71 vdd gnd cell_6t
Xbit_r72_c97 bl_97 br_97 wl_72 vdd gnd cell_6t
Xbit_r73_c97 bl_97 br_97 wl_73 vdd gnd cell_6t
Xbit_r74_c97 bl_97 br_97 wl_74 vdd gnd cell_6t
Xbit_r75_c97 bl_97 br_97 wl_75 vdd gnd cell_6t
Xbit_r76_c97 bl_97 br_97 wl_76 vdd gnd cell_6t
Xbit_r77_c97 bl_97 br_97 wl_77 vdd gnd cell_6t
Xbit_r78_c97 bl_97 br_97 wl_78 vdd gnd cell_6t
Xbit_r79_c97 bl_97 br_97 wl_79 vdd gnd cell_6t
Xbit_r80_c97 bl_97 br_97 wl_80 vdd gnd cell_6t
Xbit_r81_c97 bl_97 br_97 wl_81 vdd gnd cell_6t
Xbit_r82_c97 bl_97 br_97 wl_82 vdd gnd cell_6t
Xbit_r83_c97 bl_97 br_97 wl_83 vdd gnd cell_6t
Xbit_r84_c97 bl_97 br_97 wl_84 vdd gnd cell_6t
Xbit_r85_c97 bl_97 br_97 wl_85 vdd gnd cell_6t
Xbit_r86_c97 bl_97 br_97 wl_86 vdd gnd cell_6t
Xbit_r87_c97 bl_97 br_97 wl_87 vdd gnd cell_6t
Xbit_r88_c97 bl_97 br_97 wl_88 vdd gnd cell_6t
Xbit_r89_c97 bl_97 br_97 wl_89 vdd gnd cell_6t
Xbit_r90_c97 bl_97 br_97 wl_90 vdd gnd cell_6t
Xbit_r91_c97 bl_97 br_97 wl_91 vdd gnd cell_6t
Xbit_r92_c97 bl_97 br_97 wl_92 vdd gnd cell_6t
Xbit_r93_c97 bl_97 br_97 wl_93 vdd gnd cell_6t
Xbit_r94_c97 bl_97 br_97 wl_94 vdd gnd cell_6t
Xbit_r95_c97 bl_97 br_97 wl_95 vdd gnd cell_6t
Xbit_r96_c97 bl_97 br_97 wl_96 vdd gnd cell_6t
Xbit_r97_c97 bl_97 br_97 wl_97 vdd gnd cell_6t
Xbit_r98_c97 bl_97 br_97 wl_98 vdd gnd cell_6t
Xbit_r99_c97 bl_97 br_97 wl_99 vdd gnd cell_6t
Xbit_r100_c97 bl_97 br_97 wl_100 vdd gnd cell_6t
Xbit_r101_c97 bl_97 br_97 wl_101 vdd gnd cell_6t
Xbit_r102_c97 bl_97 br_97 wl_102 vdd gnd cell_6t
Xbit_r103_c97 bl_97 br_97 wl_103 vdd gnd cell_6t
Xbit_r104_c97 bl_97 br_97 wl_104 vdd gnd cell_6t
Xbit_r105_c97 bl_97 br_97 wl_105 vdd gnd cell_6t
Xbit_r106_c97 bl_97 br_97 wl_106 vdd gnd cell_6t
Xbit_r107_c97 bl_97 br_97 wl_107 vdd gnd cell_6t
Xbit_r108_c97 bl_97 br_97 wl_108 vdd gnd cell_6t
Xbit_r109_c97 bl_97 br_97 wl_109 vdd gnd cell_6t
Xbit_r110_c97 bl_97 br_97 wl_110 vdd gnd cell_6t
Xbit_r111_c97 bl_97 br_97 wl_111 vdd gnd cell_6t
Xbit_r112_c97 bl_97 br_97 wl_112 vdd gnd cell_6t
Xbit_r113_c97 bl_97 br_97 wl_113 vdd gnd cell_6t
Xbit_r114_c97 bl_97 br_97 wl_114 vdd gnd cell_6t
Xbit_r115_c97 bl_97 br_97 wl_115 vdd gnd cell_6t
Xbit_r116_c97 bl_97 br_97 wl_116 vdd gnd cell_6t
Xbit_r117_c97 bl_97 br_97 wl_117 vdd gnd cell_6t
Xbit_r118_c97 bl_97 br_97 wl_118 vdd gnd cell_6t
Xbit_r119_c97 bl_97 br_97 wl_119 vdd gnd cell_6t
Xbit_r120_c97 bl_97 br_97 wl_120 vdd gnd cell_6t
Xbit_r121_c97 bl_97 br_97 wl_121 vdd gnd cell_6t
Xbit_r122_c97 bl_97 br_97 wl_122 vdd gnd cell_6t
Xbit_r123_c97 bl_97 br_97 wl_123 vdd gnd cell_6t
Xbit_r124_c97 bl_97 br_97 wl_124 vdd gnd cell_6t
Xbit_r125_c97 bl_97 br_97 wl_125 vdd gnd cell_6t
Xbit_r126_c97 bl_97 br_97 wl_126 vdd gnd cell_6t
Xbit_r127_c97 bl_97 br_97 wl_127 vdd gnd cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd cell_6t
Xbit_r1_c98 bl_98 br_98 wl_1 vdd gnd cell_6t
Xbit_r2_c98 bl_98 br_98 wl_2 vdd gnd cell_6t
Xbit_r3_c98 bl_98 br_98 wl_3 vdd gnd cell_6t
Xbit_r4_c98 bl_98 br_98 wl_4 vdd gnd cell_6t
Xbit_r5_c98 bl_98 br_98 wl_5 vdd gnd cell_6t
Xbit_r6_c98 bl_98 br_98 wl_6 vdd gnd cell_6t
Xbit_r7_c98 bl_98 br_98 wl_7 vdd gnd cell_6t
Xbit_r8_c98 bl_98 br_98 wl_8 vdd gnd cell_6t
Xbit_r9_c98 bl_98 br_98 wl_9 vdd gnd cell_6t
Xbit_r10_c98 bl_98 br_98 wl_10 vdd gnd cell_6t
Xbit_r11_c98 bl_98 br_98 wl_11 vdd gnd cell_6t
Xbit_r12_c98 bl_98 br_98 wl_12 vdd gnd cell_6t
Xbit_r13_c98 bl_98 br_98 wl_13 vdd gnd cell_6t
Xbit_r14_c98 bl_98 br_98 wl_14 vdd gnd cell_6t
Xbit_r15_c98 bl_98 br_98 wl_15 vdd gnd cell_6t
Xbit_r16_c98 bl_98 br_98 wl_16 vdd gnd cell_6t
Xbit_r17_c98 bl_98 br_98 wl_17 vdd gnd cell_6t
Xbit_r18_c98 bl_98 br_98 wl_18 vdd gnd cell_6t
Xbit_r19_c98 bl_98 br_98 wl_19 vdd gnd cell_6t
Xbit_r20_c98 bl_98 br_98 wl_20 vdd gnd cell_6t
Xbit_r21_c98 bl_98 br_98 wl_21 vdd gnd cell_6t
Xbit_r22_c98 bl_98 br_98 wl_22 vdd gnd cell_6t
Xbit_r23_c98 bl_98 br_98 wl_23 vdd gnd cell_6t
Xbit_r24_c98 bl_98 br_98 wl_24 vdd gnd cell_6t
Xbit_r25_c98 bl_98 br_98 wl_25 vdd gnd cell_6t
Xbit_r26_c98 bl_98 br_98 wl_26 vdd gnd cell_6t
Xbit_r27_c98 bl_98 br_98 wl_27 vdd gnd cell_6t
Xbit_r28_c98 bl_98 br_98 wl_28 vdd gnd cell_6t
Xbit_r29_c98 bl_98 br_98 wl_29 vdd gnd cell_6t
Xbit_r30_c98 bl_98 br_98 wl_30 vdd gnd cell_6t
Xbit_r31_c98 bl_98 br_98 wl_31 vdd gnd cell_6t
Xbit_r32_c98 bl_98 br_98 wl_32 vdd gnd cell_6t
Xbit_r33_c98 bl_98 br_98 wl_33 vdd gnd cell_6t
Xbit_r34_c98 bl_98 br_98 wl_34 vdd gnd cell_6t
Xbit_r35_c98 bl_98 br_98 wl_35 vdd gnd cell_6t
Xbit_r36_c98 bl_98 br_98 wl_36 vdd gnd cell_6t
Xbit_r37_c98 bl_98 br_98 wl_37 vdd gnd cell_6t
Xbit_r38_c98 bl_98 br_98 wl_38 vdd gnd cell_6t
Xbit_r39_c98 bl_98 br_98 wl_39 vdd gnd cell_6t
Xbit_r40_c98 bl_98 br_98 wl_40 vdd gnd cell_6t
Xbit_r41_c98 bl_98 br_98 wl_41 vdd gnd cell_6t
Xbit_r42_c98 bl_98 br_98 wl_42 vdd gnd cell_6t
Xbit_r43_c98 bl_98 br_98 wl_43 vdd gnd cell_6t
Xbit_r44_c98 bl_98 br_98 wl_44 vdd gnd cell_6t
Xbit_r45_c98 bl_98 br_98 wl_45 vdd gnd cell_6t
Xbit_r46_c98 bl_98 br_98 wl_46 vdd gnd cell_6t
Xbit_r47_c98 bl_98 br_98 wl_47 vdd gnd cell_6t
Xbit_r48_c98 bl_98 br_98 wl_48 vdd gnd cell_6t
Xbit_r49_c98 bl_98 br_98 wl_49 vdd gnd cell_6t
Xbit_r50_c98 bl_98 br_98 wl_50 vdd gnd cell_6t
Xbit_r51_c98 bl_98 br_98 wl_51 vdd gnd cell_6t
Xbit_r52_c98 bl_98 br_98 wl_52 vdd gnd cell_6t
Xbit_r53_c98 bl_98 br_98 wl_53 vdd gnd cell_6t
Xbit_r54_c98 bl_98 br_98 wl_54 vdd gnd cell_6t
Xbit_r55_c98 bl_98 br_98 wl_55 vdd gnd cell_6t
Xbit_r56_c98 bl_98 br_98 wl_56 vdd gnd cell_6t
Xbit_r57_c98 bl_98 br_98 wl_57 vdd gnd cell_6t
Xbit_r58_c98 bl_98 br_98 wl_58 vdd gnd cell_6t
Xbit_r59_c98 bl_98 br_98 wl_59 vdd gnd cell_6t
Xbit_r60_c98 bl_98 br_98 wl_60 vdd gnd cell_6t
Xbit_r61_c98 bl_98 br_98 wl_61 vdd gnd cell_6t
Xbit_r62_c98 bl_98 br_98 wl_62 vdd gnd cell_6t
Xbit_r63_c98 bl_98 br_98 wl_63 vdd gnd cell_6t
Xbit_r64_c98 bl_98 br_98 wl_64 vdd gnd cell_6t
Xbit_r65_c98 bl_98 br_98 wl_65 vdd gnd cell_6t
Xbit_r66_c98 bl_98 br_98 wl_66 vdd gnd cell_6t
Xbit_r67_c98 bl_98 br_98 wl_67 vdd gnd cell_6t
Xbit_r68_c98 bl_98 br_98 wl_68 vdd gnd cell_6t
Xbit_r69_c98 bl_98 br_98 wl_69 vdd gnd cell_6t
Xbit_r70_c98 bl_98 br_98 wl_70 vdd gnd cell_6t
Xbit_r71_c98 bl_98 br_98 wl_71 vdd gnd cell_6t
Xbit_r72_c98 bl_98 br_98 wl_72 vdd gnd cell_6t
Xbit_r73_c98 bl_98 br_98 wl_73 vdd gnd cell_6t
Xbit_r74_c98 bl_98 br_98 wl_74 vdd gnd cell_6t
Xbit_r75_c98 bl_98 br_98 wl_75 vdd gnd cell_6t
Xbit_r76_c98 bl_98 br_98 wl_76 vdd gnd cell_6t
Xbit_r77_c98 bl_98 br_98 wl_77 vdd gnd cell_6t
Xbit_r78_c98 bl_98 br_98 wl_78 vdd gnd cell_6t
Xbit_r79_c98 bl_98 br_98 wl_79 vdd gnd cell_6t
Xbit_r80_c98 bl_98 br_98 wl_80 vdd gnd cell_6t
Xbit_r81_c98 bl_98 br_98 wl_81 vdd gnd cell_6t
Xbit_r82_c98 bl_98 br_98 wl_82 vdd gnd cell_6t
Xbit_r83_c98 bl_98 br_98 wl_83 vdd gnd cell_6t
Xbit_r84_c98 bl_98 br_98 wl_84 vdd gnd cell_6t
Xbit_r85_c98 bl_98 br_98 wl_85 vdd gnd cell_6t
Xbit_r86_c98 bl_98 br_98 wl_86 vdd gnd cell_6t
Xbit_r87_c98 bl_98 br_98 wl_87 vdd gnd cell_6t
Xbit_r88_c98 bl_98 br_98 wl_88 vdd gnd cell_6t
Xbit_r89_c98 bl_98 br_98 wl_89 vdd gnd cell_6t
Xbit_r90_c98 bl_98 br_98 wl_90 vdd gnd cell_6t
Xbit_r91_c98 bl_98 br_98 wl_91 vdd gnd cell_6t
Xbit_r92_c98 bl_98 br_98 wl_92 vdd gnd cell_6t
Xbit_r93_c98 bl_98 br_98 wl_93 vdd gnd cell_6t
Xbit_r94_c98 bl_98 br_98 wl_94 vdd gnd cell_6t
Xbit_r95_c98 bl_98 br_98 wl_95 vdd gnd cell_6t
Xbit_r96_c98 bl_98 br_98 wl_96 vdd gnd cell_6t
Xbit_r97_c98 bl_98 br_98 wl_97 vdd gnd cell_6t
Xbit_r98_c98 bl_98 br_98 wl_98 vdd gnd cell_6t
Xbit_r99_c98 bl_98 br_98 wl_99 vdd gnd cell_6t
Xbit_r100_c98 bl_98 br_98 wl_100 vdd gnd cell_6t
Xbit_r101_c98 bl_98 br_98 wl_101 vdd gnd cell_6t
Xbit_r102_c98 bl_98 br_98 wl_102 vdd gnd cell_6t
Xbit_r103_c98 bl_98 br_98 wl_103 vdd gnd cell_6t
Xbit_r104_c98 bl_98 br_98 wl_104 vdd gnd cell_6t
Xbit_r105_c98 bl_98 br_98 wl_105 vdd gnd cell_6t
Xbit_r106_c98 bl_98 br_98 wl_106 vdd gnd cell_6t
Xbit_r107_c98 bl_98 br_98 wl_107 vdd gnd cell_6t
Xbit_r108_c98 bl_98 br_98 wl_108 vdd gnd cell_6t
Xbit_r109_c98 bl_98 br_98 wl_109 vdd gnd cell_6t
Xbit_r110_c98 bl_98 br_98 wl_110 vdd gnd cell_6t
Xbit_r111_c98 bl_98 br_98 wl_111 vdd gnd cell_6t
Xbit_r112_c98 bl_98 br_98 wl_112 vdd gnd cell_6t
Xbit_r113_c98 bl_98 br_98 wl_113 vdd gnd cell_6t
Xbit_r114_c98 bl_98 br_98 wl_114 vdd gnd cell_6t
Xbit_r115_c98 bl_98 br_98 wl_115 vdd gnd cell_6t
Xbit_r116_c98 bl_98 br_98 wl_116 vdd gnd cell_6t
Xbit_r117_c98 bl_98 br_98 wl_117 vdd gnd cell_6t
Xbit_r118_c98 bl_98 br_98 wl_118 vdd gnd cell_6t
Xbit_r119_c98 bl_98 br_98 wl_119 vdd gnd cell_6t
Xbit_r120_c98 bl_98 br_98 wl_120 vdd gnd cell_6t
Xbit_r121_c98 bl_98 br_98 wl_121 vdd gnd cell_6t
Xbit_r122_c98 bl_98 br_98 wl_122 vdd gnd cell_6t
Xbit_r123_c98 bl_98 br_98 wl_123 vdd gnd cell_6t
Xbit_r124_c98 bl_98 br_98 wl_124 vdd gnd cell_6t
Xbit_r125_c98 bl_98 br_98 wl_125 vdd gnd cell_6t
Xbit_r126_c98 bl_98 br_98 wl_126 vdd gnd cell_6t
Xbit_r127_c98 bl_98 br_98 wl_127 vdd gnd cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd cell_6t
Xbit_r1_c99 bl_99 br_99 wl_1 vdd gnd cell_6t
Xbit_r2_c99 bl_99 br_99 wl_2 vdd gnd cell_6t
Xbit_r3_c99 bl_99 br_99 wl_3 vdd gnd cell_6t
Xbit_r4_c99 bl_99 br_99 wl_4 vdd gnd cell_6t
Xbit_r5_c99 bl_99 br_99 wl_5 vdd gnd cell_6t
Xbit_r6_c99 bl_99 br_99 wl_6 vdd gnd cell_6t
Xbit_r7_c99 bl_99 br_99 wl_7 vdd gnd cell_6t
Xbit_r8_c99 bl_99 br_99 wl_8 vdd gnd cell_6t
Xbit_r9_c99 bl_99 br_99 wl_9 vdd gnd cell_6t
Xbit_r10_c99 bl_99 br_99 wl_10 vdd gnd cell_6t
Xbit_r11_c99 bl_99 br_99 wl_11 vdd gnd cell_6t
Xbit_r12_c99 bl_99 br_99 wl_12 vdd gnd cell_6t
Xbit_r13_c99 bl_99 br_99 wl_13 vdd gnd cell_6t
Xbit_r14_c99 bl_99 br_99 wl_14 vdd gnd cell_6t
Xbit_r15_c99 bl_99 br_99 wl_15 vdd gnd cell_6t
Xbit_r16_c99 bl_99 br_99 wl_16 vdd gnd cell_6t
Xbit_r17_c99 bl_99 br_99 wl_17 vdd gnd cell_6t
Xbit_r18_c99 bl_99 br_99 wl_18 vdd gnd cell_6t
Xbit_r19_c99 bl_99 br_99 wl_19 vdd gnd cell_6t
Xbit_r20_c99 bl_99 br_99 wl_20 vdd gnd cell_6t
Xbit_r21_c99 bl_99 br_99 wl_21 vdd gnd cell_6t
Xbit_r22_c99 bl_99 br_99 wl_22 vdd gnd cell_6t
Xbit_r23_c99 bl_99 br_99 wl_23 vdd gnd cell_6t
Xbit_r24_c99 bl_99 br_99 wl_24 vdd gnd cell_6t
Xbit_r25_c99 bl_99 br_99 wl_25 vdd gnd cell_6t
Xbit_r26_c99 bl_99 br_99 wl_26 vdd gnd cell_6t
Xbit_r27_c99 bl_99 br_99 wl_27 vdd gnd cell_6t
Xbit_r28_c99 bl_99 br_99 wl_28 vdd gnd cell_6t
Xbit_r29_c99 bl_99 br_99 wl_29 vdd gnd cell_6t
Xbit_r30_c99 bl_99 br_99 wl_30 vdd gnd cell_6t
Xbit_r31_c99 bl_99 br_99 wl_31 vdd gnd cell_6t
Xbit_r32_c99 bl_99 br_99 wl_32 vdd gnd cell_6t
Xbit_r33_c99 bl_99 br_99 wl_33 vdd gnd cell_6t
Xbit_r34_c99 bl_99 br_99 wl_34 vdd gnd cell_6t
Xbit_r35_c99 bl_99 br_99 wl_35 vdd gnd cell_6t
Xbit_r36_c99 bl_99 br_99 wl_36 vdd gnd cell_6t
Xbit_r37_c99 bl_99 br_99 wl_37 vdd gnd cell_6t
Xbit_r38_c99 bl_99 br_99 wl_38 vdd gnd cell_6t
Xbit_r39_c99 bl_99 br_99 wl_39 vdd gnd cell_6t
Xbit_r40_c99 bl_99 br_99 wl_40 vdd gnd cell_6t
Xbit_r41_c99 bl_99 br_99 wl_41 vdd gnd cell_6t
Xbit_r42_c99 bl_99 br_99 wl_42 vdd gnd cell_6t
Xbit_r43_c99 bl_99 br_99 wl_43 vdd gnd cell_6t
Xbit_r44_c99 bl_99 br_99 wl_44 vdd gnd cell_6t
Xbit_r45_c99 bl_99 br_99 wl_45 vdd gnd cell_6t
Xbit_r46_c99 bl_99 br_99 wl_46 vdd gnd cell_6t
Xbit_r47_c99 bl_99 br_99 wl_47 vdd gnd cell_6t
Xbit_r48_c99 bl_99 br_99 wl_48 vdd gnd cell_6t
Xbit_r49_c99 bl_99 br_99 wl_49 vdd gnd cell_6t
Xbit_r50_c99 bl_99 br_99 wl_50 vdd gnd cell_6t
Xbit_r51_c99 bl_99 br_99 wl_51 vdd gnd cell_6t
Xbit_r52_c99 bl_99 br_99 wl_52 vdd gnd cell_6t
Xbit_r53_c99 bl_99 br_99 wl_53 vdd gnd cell_6t
Xbit_r54_c99 bl_99 br_99 wl_54 vdd gnd cell_6t
Xbit_r55_c99 bl_99 br_99 wl_55 vdd gnd cell_6t
Xbit_r56_c99 bl_99 br_99 wl_56 vdd gnd cell_6t
Xbit_r57_c99 bl_99 br_99 wl_57 vdd gnd cell_6t
Xbit_r58_c99 bl_99 br_99 wl_58 vdd gnd cell_6t
Xbit_r59_c99 bl_99 br_99 wl_59 vdd gnd cell_6t
Xbit_r60_c99 bl_99 br_99 wl_60 vdd gnd cell_6t
Xbit_r61_c99 bl_99 br_99 wl_61 vdd gnd cell_6t
Xbit_r62_c99 bl_99 br_99 wl_62 vdd gnd cell_6t
Xbit_r63_c99 bl_99 br_99 wl_63 vdd gnd cell_6t
Xbit_r64_c99 bl_99 br_99 wl_64 vdd gnd cell_6t
Xbit_r65_c99 bl_99 br_99 wl_65 vdd gnd cell_6t
Xbit_r66_c99 bl_99 br_99 wl_66 vdd gnd cell_6t
Xbit_r67_c99 bl_99 br_99 wl_67 vdd gnd cell_6t
Xbit_r68_c99 bl_99 br_99 wl_68 vdd gnd cell_6t
Xbit_r69_c99 bl_99 br_99 wl_69 vdd gnd cell_6t
Xbit_r70_c99 bl_99 br_99 wl_70 vdd gnd cell_6t
Xbit_r71_c99 bl_99 br_99 wl_71 vdd gnd cell_6t
Xbit_r72_c99 bl_99 br_99 wl_72 vdd gnd cell_6t
Xbit_r73_c99 bl_99 br_99 wl_73 vdd gnd cell_6t
Xbit_r74_c99 bl_99 br_99 wl_74 vdd gnd cell_6t
Xbit_r75_c99 bl_99 br_99 wl_75 vdd gnd cell_6t
Xbit_r76_c99 bl_99 br_99 wl_76 vdd gnd cell_6t
Xbit_r77_c99 bl_99 br_99 wl_77 vdd gnd cell_6t
Xbit_r78_c99 bl_99 br_99 wl_78 vdd gnd cell_6t
Xbit_r79_c99 bl_99 br_99 wl_79 vdd gnd cell_6t
Xbit_r80_c99 bl_99 br_99 wl_80 vdd gnd cell_6t
Xbit_r81_c99 bl_99 br_99 wl_81 vdd gnd cell_6t
Xbit_r82_c99 bl_99 br_99 wl_82 vdd gnd cell_6t
Xbit_r83_c99 bl_99 br_99 wl_83 vdd gnd cell_6t
Xbit_r84_c99 bl_99 br_99 wl_84 vdd gnd cell_6t
Xbit_r85_c99 bl_99 br_99 wl_85 vdd gnd cell_6t
Xbit_r86_c99 bl_99 br_99 wl_86 vdd gnd cell_6t
Xbit_r87_c99 bl_99 br_99 wl_87 vdd gnd cell_6t
Xbit_r88_c99 bl_99 br_99 wl_88 vdd gnd cell_6t
Xbit_r89_c99 bl_99 br_99 wl_89 vdd gnd cell_6t
Xbit_r90_c99 bl_99 br_99 wl_90 vdd gnd cell_6t
Xbit_r91_c99 bl_99 br_99 wl_91 vdd gnd cell_6t
Xbit_r92_c99 bl_99 br_99 wl_92 vdd gnd cell_6t
Xbit_r93_c99 bl_99 br_99 wl_93 vdd gnd cell_6t
Xbit_r94_c99 bl_99 br_99 wl_94 vdd gnd cell_6t
Xbit_r95_c99 bl_99 br_99 wl_95 vdd gnd cell_6t
Xbit_r96_c99 bl_99 br_99 wl_96 vdd gnd cell_6t
Xbit_r97_c99 bl_99 br_99 wl_97 vdd gnd cell_6t
Xbit_r98_c99 bl_99 br_99 wl_98 vdd gnd cell_6t
Xbit_r99_c99 bl_99 br_99 wl_99 vdd gnd cell_6t
Xbit_r100_c99 bl_99 br_99 wl_100 vdd gnd cell_6t
Xbit_r101_c99 bl_99 br_99 wl_101 vdd gnd cell_6t
Xbit_r102_c99 bl_99 br_99 wl_102 vdd gnd cell_6t
Xbit_r103_c99 bl_99 br_99 wl_103 vdd gnd cell_6t
Xbit_r104_c99 bl_99 br_99 wl_104 vdd gnd cell_6t
Xbit_r105_c99 bl_99 br_99 wl_105 vdd gnd cell_6t
Xbit_r106_c99 bl_99 br_99 wl_106 vdd gnd cell_6t
Xbit_r107_c99 bl_99 br_99 wl_107 vdd gnd cell_6t
Xbit_r108_c99 bl_99 br_99 wl_108 vdd gnd cell_6t
Xbit_r109_c99 bl_99 br_99 wl_109 vdd gnd cell_6t
Xbit_r110_c99 bl_99 br_99 wl_110 vdd gnd cell_6t
Xbit_r111_c99 bl_99 br_99 wl_111 vdd gnd cell_6t
Xbit_r112_c99 bl_99 br_99 wl_112 vdd gnd cell_6t
Xbit_r113_c99 bl_99 br_99 wl_113 vdd gnd cell_6t
Xbit_r114_c99 bl_99 br_99 wl_114 vdd gnd cell_6t
Xbit_r115_c99 bl_99 br_99 wl_115 vdd gnd cell_6t
Xbit_r116_c99 bl_99 br_99 wl_116 vdd gnd cell_6t
Xbit_r117_c99 bl_99 br_99 wl_117 vdd gnd cell_6t
Xbit_r118_c99 bl_99 br_99 wl_118 vdd gnd cell_6t
Xbit_r119_c99 bl_99 br_99 wl_119 vdd gnd cell_6t
Xbit_r120_c99 bl_99 br_99 wl_120 vdd gnd cell_6t
Xbit_r121_c99 bl_99 br_99 wl_121 vdd gnd cell_6t
Xbit_r122_c99 bl_99 br_99 wl_122 vdd gnd cell_6t
Xbit_r123_c99 bl_99 br_99 wl_123 vdd gnd cell_6t
Xbit_r124_c99 bl_99 br_99 wl_124 vdd gnd cell_6t
Xbit_r125_c99 bl_99 br_99 wl_125 vdd gnd cell_6t
Xbit_r126_c99 bl_99 br_99 wl_126 vdd gnd cell_6t
Xbit_r127_c99 bl_99 br_99 wl_127 vdd gnd cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd cell_6t
Xbit_r1_c100 bl_100 br_100 wl_1 vdd gnd cell_6t
Xbit_r2_c100 bl_100 br_100 wl_2 vdd gnd cell_6t
Xbit_r3_c100 bl_100 br_100 wl_3 vdd gnd cell_6t
Xbit_r4_c100 bl_100 br_100 wl_4 vdd gnd cell_6t
Xbit_r5_c100 bl_100 br_100 wl_5 vdd gnd cell_6t
Xbit_r6_c100 bl_100 br_100 wl_6 vdd gnd cell_6t
Xbit_r7_c100 bl_100 br_100 wl_7 vdd gnd cell_6t
Xbit_r8_c100 bl_100 br_100 wl_8 vdd gnd cell_6t
Xbit_r9_c100 bl_100 br_100 wl_9 vdd gnd cell_6t
Xbit_r10_c100 bl_100 br_100 wl_10 vdd gnd cell_6t
Xbit_r11_c100 bl_100 br_100 wl_11 vdd gnd cell_6t
Xbit_r12_c100 bl_100 br_100 wl_12 vdd gnd cell_6t
Xbit_r13_c100 bl_100 br_100 wl_13 vdd gnd cell_6t
Xbit_r14_c100 bl_100 br_100 wl_14 vdd gnd cell_6t
Xbit_r15_c100 bl_100 br_100 wl_15 vdd gnd cell_6t
Xbit_r16_c100 bl_100 br_100 wl_16 vdd gnd cell_6t
Xbit_r17_c100 bl_100 br_100 wl_17 vdd gnd cell_6t
Xbit_r18_c100 bl_100 br_100 wl_18 vdd gnd cell_6t
Xbit_r19_c100 bl_100 br_100 wl_19 vdd gnd cell_6t
Xbit_r20_c100 bl_100 br_100 wl_20 vdd gnd cell_6t
Xbit_r21_c100 bl_100 br_100 wl_21 vdd gnd cell_6t
Xbit_r22_c100 bl_100 br_100 wl_22 vdd gnd cell_6t
Xbit_r23_c100 bl_100 br_100 wl_23 vdd gnd cell_6t
Xbit_r24_c100 bl_100 br_100 wl_24 vdd gnd cell_6t
Xbit_r25_c100 bl_100 br_100 wl_25 vdd gnd cell_6t
Xbit_r26_c100 bl_100 br_100 wl_26 vdd gnd cell_6t
Xbit_r27_c100 bl_100 br_100 wl_27 vdd gnd cell_6t
Xbit_r28_c100 bl_100 br_100 wl_28 vdd gnd cell_6t
Xbit_r29_c100 bl_100 br_100 wl_29 vdd gnd cell_6t
Xbit_r30_c100 bl_100 br_100 wl_30 vdd gnd cell_6t
Xbit_r31_c100 bl_100 br_100 wl_31 vdd gnd cell_6t
Xbit_r32_c100 bl_100 br_100 wl_32 vdd gnd cell_6t
Xbit_r33_c100 bl_100 br_100 wl_33 vdd gnd cell_6t
Xbit_r34_c100 bl_100 br_100 wl_34 vdd gnd cell_6t
Xbit_r35_c100 bl_100 br_100 wl_35 vdd gnd cell_6t
Xbit_r36_c100 bl_100 br_100 wl_36 vdd gnd cell_6t
Xbit_r37_c100 bl_100 br_100 wl_37 vdd gnd cell_6t
Xbit_r38_c100 bl_100 br_100 wl_38 vdd gnd cell_6t
Xbit_r39_c100 bl_100 br_100 wl_39 vdd gnd cell_6t
Xbit_r40_c100 bl_100 br_100 wl_40 vdd gnd cell_6t
Xbit_r41_c100 bl_100 br_100 wl_41 vdd gnd cell_6t
Xbit_r42_c100 bl_100 br_100 wl_42 vdd gnd cell_6t
Xbit_r43_c100 bl_100 br_100 wl_43 vdd gnd cell_6t
Xbit_r44_c100 bl_100 br_100 wl_44 vdd gnd cell_6t
Xbit_r45_c100 bl_100 br_100 wl_45 vdd gnd cell_6t
Xbit_r46_c100 bl_100 br_100 wl_46 vdd gnd cell_6t
Xbit_r47_c100 bl_100 br_100 wl_47 vdd gnd cell_6t
Xbit_r48_c100 bl_100 br_100 wl_48 vdd gnd cell_6t
Xbit_r49_c100 bl_100 br_100 wl_49 vdd gnd cell_6t
Xbit_r50_c100 bl_100 br_100 wl_50 vdd gnd cell_6t
Xbit_r51_c100 bl_100 br_100 wl_51 vdd gnd cell_6t
Xbit_r52_c100 bl_100 br_100 wl_52 vdd gnd cell_6t
Xbit_r53_c100 bl_100 br_100 wl_53 vdd gnd cell_6t
Xbit_r54_c100 bl_100 br_100 wl_54 vdd gnd cell_6t
Xbit_r55_c100 bl_100 br_100 wl_55 vdd gnd cell_6t
Xbit_r56_c100 bl_100 br_100 wl_56 vdd gnd cell_6t
Xbit_r57_c100 bl_100 br_100 wl_57 vdd gnd cell_6t
Xbit_r58_c100 bl_100 br_100 wl_58 vdd gnd cell_6t
Xbit_r59_c100 bl_100 br_100 wl_59 vdd gnd cell_6t
Xbit_r60_c100 bl_100 br_100 wl_60 vdd gnd cell_6t
Xbit_r61_c100 bl_100 br_100 wl_61 vdd gnd cell_6t
Xbit_r62_c100 bl_100 br_100 wl_62 vdd gnd cell_6t
Xbit_r63_c100 bl_100 br_100 wl_63 vdd gnd cell_6t
Xbit_r64_c100 bl_100 br_100 wl_64 vdd gnd cell_6t
Xbit_r65_c100 bl_100 br_100 wl_65 vdd gnd cell_6t
Xbit_r66_c100 bl_100 br_100 wl_66 vdd gnd cell_6t
Xbit_r67_c100 bl_100 br_100 wl_67 vdd gnd cell_6t
Xbit_r68_c100 bl_100 br_100 wl_68 vdd gnd cell_6t
Xbit_r69_c100 bl_100 br_100 wl_69 vdd gnd cell_6t
Xbit_r70_c100 bl_100 br_100 wl_70 vdd gnd cell_6t
Xbit_r71_c100 bl_100 br_100 wl_71 vdd gnd cell_6t
Xbit_r72_c100 bl_100 br_100 wl_72 vdd gnd cell_6t
Xbit_r73_c100 bl_100 br_100 wl_73 vdd gnd cell_6t
Xbit_r74_c100 bl_100 br_100 wl_74 vdd gnd cell_6t
Xbit_r75_c100 bl_100 br_100 wl_75 vdd gnd cell_6t
Xbit_r76_c100 bl_100 br_100 wl_76 vdd gnd cell_6t
Xbit_r77_c100 bl_100 br_100 wl_77 vdd gnd cell_6t
Xbit_r78_c100 bl_100 br_100 wl_78 vdd gnd cell_6t
Xbit_r79_c100 bl_100 br_100 wl_79 vdd gnd cell_6t
Xbit_r80_c100 bl_100 br_100 wl_80 vdd gnd cell_6t
Xbit_r81_c100 bl_100 br_100 wl_81 vdd gnd cell_6t
Xbit_r82_c100 bl_100 br_100 wl_82 vdd gnd cell_6t
Xbit_r83_c100 bl_100 br_100 wl_83 vdd gnd cell_6t
Xbit_r84_c100 bl_100 br_100 wl_84 vdd gnd cell_6t
Xbit_r85_c100 bl_100 br_100 wl_85 vdd gnd cell_6t
Xbit_r86_c100 bl_100 br_100 wl_86 vdd gnd cell_6t
Xbit_r87_c100 bl_100 br_100 wl_87 vdd gnd cell_6t
Xbit_r88_c100 bl_100 br_100 wl_88 vdd gnd cell_6t
Xbit_r89_c100 bl_100 br_100 wl_89 vdd gnd cell_6t
Xbit_r90_c100 bl_100 br_100 wl_90 vdd gnd cell_6t
Xbit_r91_c100 bl_100 br_100 wl_91 vdd gnd cell_6t
Xbit_r92_c100 bl_100 br_100 wl_92 vdd gnd cell_6t
Xbit_r93_c100 bl_100 br_100 wl_93 vdd gnd cell_6t
Xbit_r94_c100 bl_100 br_100 wl_94 vdd gnd cell_6t
Xbit_r95_c100 bl_100 br_100 wl_95 vdd gnd cell_6t
Xbit_r96_c100 bl_100 br_100 wl_96 vdd gnd cell_6t
Xbit_r97_c100 bl_100 br_100 wl_97 vdd gnd cell_6t
Xbit_r98_c100 bl_100 br_100 wl_98 vdd gnd cell_6t
Xbit_r99_c100 bl_100 br_100 wl_99 vdd gnd cell_6t
Xbit_r100_c100 bl_100 br_100 wl_100 vdd gnd cell_6t
Xbit_r101_c100 bl_100 br_100 wl_101 vdd gnd cell_6t
Xbit_r102_c100 bl_100 br_100 wl_102 vdd gnd cell_6t
Xbit_r103_c100 bl_100 br_100 wl_103 vdd gnd cell_6t
Xbit_r104_c100 bl_100 br_100 wl_104 vdd gnd cell_6t
Xbit_r105_c100 bl_100 br_100 wl_105 vdd gnd cell_6t
Xbit_r106_c100 bl_100 br_100 wl_106 vdd gnd cell_6t
Xbit_r107_c100 bl_100 br_100 wl_107 vdd gnd cell_6t
Xbit_r108_c100 bl_100 br_100 wl_108 vdd gnd cell_6t
Xbit_r109_c100 bl_100 br_100 wl_109 vdd gnd cell_6t
Xbit_r110_c100 bl_100 br_100 wl_110 vdd gnd cell_6t
Xbit_r111_c100 bl_100 br_100 wl_111 vdd gnd cell_6t
Xbit_r112_c100 bl_100 br_100 wl_112 vdd gnd cell_6t
Xbit_r113_c100 bl_100 br_100 wl_113 vdd gnd cell_6t
Xbit_r114_c100 bl_100 br_100 wl_114 vdd gnd cell_6t
Xbit_r115_c100 bl_100 br_100 wl_115 vdd gnd cell_6t
Xbit_r116_c100 bl_100 br_100 wl_116 vdd gnd cell_6t
Xbit_r117_c100 bl_100 br_100 wl_117 vdd gnd cell_6t
Xbit_r118_c100 bl_100 br_100 wl_118 vdd gnd cell_6t
Xbit_r119_c100 bl_100 br_100 wl_119 vdd gnd cell_6t
Xbit_r120_c100 bl_100 br_100 wl_120 vdd gnd cell_6t
Xbit_r121_c100 bl_100 br_100 wl_121 vdd gnd cell_6t
Xbit_r122_c100 bl_100 br_100 wl_122 vdd gnd cell_6t
Xbit_r123_c100 bl_100 br_100 wl_123 vdd gnd cell_6t
Xbit_r124_c100 bl_100 br_100 wl_124 vdd gnd cell_6t
Xbit_r125_c100 bl_100 br_100 wl_125 vdd gnd cell_6t
Xbit_r126_c100 bl_100 br_100 wl_126 vdd gnd cell_6t
Xbit_r127_c100 bl_100 br_100 wl_127 vdd gnd cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd cell_6t
Xbit_r1_c101 bl_101 br_101 wl_1 vdd gnd cell_6t
Xbit_r2_c101 bl_101 br_101 wl_2 vdd gnd cell_6t
Xbit_r3_c101 bl_101 br_101 wl_3 vdd gnd cell_6t
Xbit_r4_c101 bl_101 br_101 wl_4 vdd gnd cell_6t
Xbit_r5_c101 bl_101 br_101 wl_5 vdd gnd cell_6t
Xbit_r6_c101 bl_101 br_101 wl_6 vdd gnd cell_6t
Xbit_r7_c101 bl_101 br_101 wl_7 vdd gnd cell_6t
Xbit_r8_c101 bl_101 br_101 wl_8 vdd gnd cell_6t
Xbit_r9_c101 bl_101 br_101 wl_9 vdd gnd cell_6t
Xbit_r10_c101 bl_101 br_101 wl_10 vdd gnd cell_6t
Xbit_r11_c101 bl_101 br_101 wl_11 vdd gnd cell_6t
Xbit_r12_c101 bl_101 br_101 wl_12 vdd gnd cell_6t
Xbit_r13_c101 bl_101 br_101 wl_13 vdd gnd cell_6t
Xbit_r14_c101 bl_101 br_101 wl_14 vdd gnd cell_6t
Xbit_r15_c101 bl_101 br_101 wl_15 vdd gnd cell_6t
Xbit_r16_c101 bl_101 br_101 wl_16 vdd gnd cell_6t
Xbit_r17_c101 bl_101 br_101 wl_17 vdd gnd cell_6t
Xbit_r18_c101 bl_101 br_101 wl_18 vdd gnd cell_6t
Xbit_r19_c101 bl_101 br_101 wl_19 vdd gnd cell_6t
Xbit_r20_c101 bl_101 br_101 wl_20 vdd gnd cell_6t
Xbit_r21_c101 bl_101 br_101 wl_21 vdd gnd cell_6t
Xbit_r22_c101 bl_101 br_101 wl_22 vdd gnd cell_6t
Xbit_r23_c101 bl_101 br_101 wl_23 vdd gnd cell_6t
Xbit_r24_c101 bl_101 br_101 wl_24 vdd gnd cell_6t
Xbit_r25_c101 bl_101 br_101 wl_25 vdd gnd cell_6t
Xbit_r26_c101 bl_101 br_101 wl_26 vdd gnd cell_6t
Xbit_r27_c101 bl_101 br_101 wl_27 vdd gnd cell_6t
Xbit_r28_c101 bl_101 br_101 wl_28 vdd gnd cell_6t
Xbit_r29_c101 bl_101 br_101 wl_29 vdd gnd cell_6t
Xbit_r30_c101 bl_101 br_101 wl_30 vdd gnd cell_6t
Xbit_r31_c101 bl_101 br_101 wl_31 vdd gnd cell_6t
Xbit_r32_c101 bl_101 br_101 wl_32 vdd gnd cell_6t
Xbit_r33_c101 bl_101 br_101 wl_33 vdd gnd cell_6t
Xbit_r34_c101 bl_101 br_101 wl_34 vdd gnd cell_6t
Xbit_r35_c101 bl_101 br_101 wl_35 vdd gnd cell_6t
Xbit_r36_c101 bl_101 br_101 wl_36 vdd gnd cell_6t
Xbit_r37_c101 bl_101 br_101 wl_37 vdd gnd cell_6t
Xbit_r38_c101 bl_101 br_101 wl_38 vdd gnd cell_6t
Xbit_r39_c101 bl_101 br_101 wl_39 vdd gnd cell_6t
Xbit_r40_c101 bl_101 br_101 wl_40 vdd gnd cell_6t
Xbit_r41_c101 bl_101 br_101 wl_41 vdd gnd cell_6t
Xbit_r42_c101 bl_101 br_101 wl_42 vdd gnd cell_6t
Xbit_r43_c101 bl_101 br_101 wl_43 vdd gnd cell_6t
Xbit_r44_c101 bl_101 br_101 wl_44 vdd gnd cell_6t
Xbit_r45_c101 bl_101 br_101 wl_45 vdd gnd cell_6t
Xbit_r46_c101 bl_101 br_101 wl_46 vdd gnd cell_6t
Xbit_r47_c101 bl_101 br_101 wl_47 vdd gnd cell_6t
Xbit_r48_c101 bl_101 br_101 wl_48 vdd gnd cell_6t
Xbit_r49_c101 bl_101 br_101 wl_49 vdd gnd cell_6t
Xbit_r50_c101 bl_101 br_101 wl_50 vdd gnd cell_6t
Xbit_r51_c101 bl_101 br_101 wl_51 vdd gnd cell_6t
Xbit_r52_c101 bl_101 br_101 wl_52 vdd gnd cell_6t
Xbit_r53_c101 bl_101 br_101 wl_53 vdd gnd cell_6t
Xbit_r54_c101 bl_101 br_101 wl_54 vdd gnd cell_6t
Xbit_r55_c101 bl_101 br_101 wl_55 vdd gnd cell_6t
Xbit_r56_c101 bl_101 br_101 wl_56 vdd gnd cell_6t
Xbit_r57_c101 bl_101 br_101 wl_57 vdd gnd cell_6t
Xbit_r58_c101 bl_101 br_101 wl_58 vdd gnd cell_6t
Xbit_r59_c101 bl_101 br_101 wl_59 vdd gnd cell_6t
Xbit_r60_c101 bl_101 br_101 wl_60 vdd gnd cell_6t
Xbit_r61_c101 bl_101 br_101 wl_61 vdd gnd cell_6t
Xbit_r62_c101 bl_101 br_101 wl_62 vdd gnd cell_6t
Xbit_r63_c101 bl_101 br_101 wl_63 vdd gnd cell_6t
Xbit_r64_c101 bl_101 br_101 wl_64 vdd gnd cell_6t
Xbit_r65_c101 bl_101 br_101 wl_65 vdd gnd cell_6t
Xbit_r66_c101 bl_101 br_101 wl_66 vdd gnd cell_6t
Xbit_r67_c101 bl_101 br_101 wl_67 vdd gnd cell_6t
Xbit_r68_c101 bl_101 br_101 wl_68 vdd gnd cell_6t
Xbit_r69_c101 bl_101 br_101 wl_69 vdd gnd cell_6t
Xbit_r70_c101 bl_101 br_101 wl_70 vdd gnd cell_6t
Xbit_r71_c101 bl_101 br_101 wl_71 vdd gnd cell_6t
Xbit_r72_c101 bl_101 br_101 wl_72 vdd gnd cell_6t
Xbit_r73_c101 bl_101 br_101 wl_73 vdd gnd cell_6t
Xbit_r74_c101 bl_101 br_101 wl_74 vdd gnd cell_6t
Xbit_r75_c101 bl_101 br_101 wl_75 vdd gnd cell_6t
Xbit_r76_c101 bl_101 br_101 wl_76 vdd gnd cell_6t
Xbit_r77_c101 bl_101 br_101 wl_77 vdd gnd cell_6t
Xbit_r78_c101 bl_101 br_101 wl_78 vdd gnd cell_6t
Xbit_r79_c101 bl_101 br_101 wl_79 vdd gnd cell_6t
Xbit_r80_c101 bl_101 br_101 wl_80 vdd gnd cell_6t
Xbit_r81_c101 bl_101 br_101 wl_81 vdd gnd cell_6t
Xbit_r82_c101 bl_101 br_101 wl_82 vdd gnd cell_6t
Xbit_r83_c101 bl_101 br_101 wl_83 vdd gnd cell_6t
Xbit_r84_c101 bl_101 br_101 wl_84 vdd gnd cell_6t
Xbit_r85_c101 bl_101 br_101 wl_85 vdd gnd cell_6t
Xbit_r86_c101 bl_101 br_101 wl_86 vdd gnd cell_6t
Xbit_r87_c101 bl_101 br_101 wl_87 vdd gnd cell_6t
Xbit_r88_c101 bl_101 br_101 wl_88 vdd gnd cell_6t
Xbit_r89_c101 bl_101 br_101 wl_89 vdd gnd cell_6t
Xbit_r90_c101 bl_101 br_101 wl_90 vdd gnd cell_6t
Xbit_r91_c101 bl_101 br_101 wl_91 vdd gnd cell_6t
Xbit_r92_c101 bl_101 br_101 wl_92 vdd gnd cell_6t
Xbit_r93_c101 bl_101 br_101 wl_93 vdd gnd cell_6t
Xbit_r94_c101 bl_101 br_101 wl_94 vdd gnd cell_6t
Xbit_r95_c101 bl_101 br_101 wl_95 vdd gnd cell_6t
Xbit_r96_c101 bl_101 br_101 wl_96 vdd gnd cell_6t
Xbit_r97_c101 bl_101 br_101 wl_97 vdd gnd cell_6t
Xbit_r98_c101 bl_101 br_101 wl_98 vdd gnd cell_6t
Xbit_r99_c101 bl_101 br_101 wl_99 vdd gnd cell_6t
Xbit_r100_c101 bl_101 br_101 wl_100 vdd gnd cell_6t
Xbit_r101_c101 bl_101 br_101 wl_101 vdd gnd cell_6t
Xbit_r102_c101 bl_101 br_101 wl_102 vdd gnd cell_6t
Xbit_r103_c101 bl_101 br_101 wl_103 vdd gnd cell_6t
Xbit_r104_c101 bl_101 br_101 wl_104 vdd gnd cell_6t
Xbit_r105_c101 bl_101 br_101 wl_105 vdd gnd cell_6t
Xbit_r106_c101 bl_101 br_101 wl_106 vdd gnd cell_6t
Xbit_r107_c101 bl_101 br_101 wl_107 vdd gnd cell_6t
Xbit_r108_c101 bl_101 br_101 wl_108 vdd gnd cell_6t
Xbit_r109_c101 bl_101 br_101 wl_109 vdd gnd cell_6t
Xbit_r110_c101 bl_101 br_101 wl_110 vdd gnd cell_6t
Xbit_r111_c101 bl_101 br_101 wl_111 vdd gnd cell_6t
Xbit_r112_c101 bl_101 br_101 wl_112 vdd gnd cell_6t
Xbit_r113_c101 bl_101 br_101 wl_113 vdd gnd cell_6t
Xbit_r114_c101 bl_101 br_101 wl_114 vdd gnd cell_6t
Xbit_r115_c101 bl_101 br_101 wl_115 vdd gnd cell_6t
Xbit_r116_c101 bl_101 br_101 wl_116 vdd gnd cell_6t
Xbit_r117_c101 bl_101 br_101 wl_117 vdd gnd cell_6t
Xbit_r118_c101 bl_101 br_101 wl_118 vdd gnd cell_6t
Xbit_r119_c101 bl_101 br_101 wl_119 vdd gnd cell_6t
Xbit_r120_c101 bl_101 br_101 wl_120 vdd gnd cell_6t
Xbit_r121_c101 bl_101 br_101 wl_121 vdd gnd cell_6t
Xbit_r122_c101 bl_101 br_101 wl_122 vdd gnd cell_6t
Xbit_r123_c101 bl_101 br_101 wl_123 vdd gnd cell_6t
Xbit_r124_c101 bl_101 br_101 wl_124 vdd gnd cell_6t
Xbit_r125_c101 bl_101 br_101 wl_125 vdd gnd cell_6t
Xbit_r126_c101 bl_101 br_101 wl_126 vdd gnd cell_6t
Xbit_r127_c101 bl_101 br_101 wl_127 vdd gnd cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd cell_6t
Xbit_r1_c102 bl_102 br_102 wl_1 vdd gnd cell_6t
Xbit_r2_c102 bl_102 br_102 wl_2 vdd gnd cell_6t
Xbit_r3_c102 bl_102 br_102 wl_3 vdd gnd cell_6t
Xbit_r4_c102 bl_102 br_102 wl_4 vdd gnd cell_6t
Xbit_r5_c102 bl_102 br_102 wl_5 vdd gnd cell_6t
Xbit_r6_c102 bl_102 br_102 wl_6 vdd gnd cell_6t
Xbit_r7_c102 bl_102 br_102 wl_7 vdd gnd cell_6t
Xbit_r8_c102 bl_102 br_102 wl_8 vdd gnd cell_6t
Xbit_r9_c102 bl_102 br_102 wl_9 vdd gnd cell_6t
Xbit_r10_c102 bl_102 br_102 wl_10 vdd gnd cell_6t
Xbit_r11_c102 bl_102 br_102 wl_11 vdd gnd cell_6t
Xbit_r12_c102 bl_102 br_102 wl_12 vdd gnd cell_6t
Xbit_r13_c102 bl_102 br_102 wl_13 vdd gnd cell_6t
Xbit_r14_c102 bl_102 br_102 wl_14 vdd gnd cell_6t
Xbit_r15_c102 bl_102 br_102 wl_15 vdd gnd cell_6t
Xbit_r16_c102 bl_102 br_102 wl_16 vdd gnd cell_6t
Xbit_r17_c102 bl_102 br_102 wl_17 vdd gnd cell_6t
Xbit_r18_c102 bl_102 br_102 wl_18 vdd gnd cell_6t
Xbit_r19_c102 bl_102 br_102 wl_19 vdd gnd cell_6t
Xbit_r20_c102 bl_102 br_102 wl_20 vdd gnd cell_6t
Xbit_r21_c102 bl_102 br_102 wl_21 vdd gnd cell_6t
Xbit_r22_c102 bl_102 br_102 wl_22 vdd gnd cell_6t
Xbit_r23_c102 bl_102 br_102 wl_23 vdd gnd cell_6t
Xbit_r24_c102 bl_102 br_102 wl_24 vdd gnd cell_6t
Xbit_r25_c102 bl_102 br_102 wl_25 vdd gnd cell_6t
Xbit_r26_c102 bl_102 br_102 wl_26 vdd gnd cell_6t
Xbit_r27_c102 bl_102 br_102 wl_27 vdd gnd cell_6t
Xbit_r28_c102 bl_102 br_102 wl_28 vdd gnd cell_6t
Xbit_r29_c102 bl_102 br_102 wl_29 vdd gnd cell_6t
Xbit_r30_c102 bl_102 br_102 wl_30 vdd gnd cell_6t
Xbit_r31_c102 bl_102 br_102 wl_31 vdd gnd cell_6t
Xbit_r32_c102 bl_102 br_102 wl_32 vdd gnd cell_6t
Xbit_r33_c102 bl_102 br_102 wl_33 vdd gnd cell_6t
Xbit_r34_c102 bl_102 br_102 wl_34 vdd gnd cell_6t
Xbit_r35_c102 bl_102 br_102 wl_35 vdd gnd cell_6t
Xbit_r36_c102 bl_102 br_102 wl_36 vdd gnd cell_6t
Xbit_r37_c102 bl_102 br_102 wl_37 vdd gnd cell_6t
Xbit_r38_c102 bl_102 br_102 wl_38 vdd gnd cell_6t
Xbit_r39_c102 bl_102 br_102 wl_39 vdd gnd cell_6t
Xbit_r40_c102 bl_102 br_102 wl_40 vdd gnd cell_6t
Xbit_r41_c102 bl_102 br_102 wl_41 vdd gnd cell_6t
Xbit_r42_c102 bl_102 br_102 wl_42 vdd gnd cell_6t
Xbit_r43_c102 bl_102 br_102 wl_43 vdd gnd cell_6t
Xbit_r44_c102 bl_102 br_102 wl_44 vdd gnd cell_6t
Xbit_r45_c102 bl_102 br_102 wl_45 vdd gnd cell_6t
Xbit_r46_c102 bl_102 br_102 wl_46 vdd gnd cell_6t
Xbit_r47_c102 bl_102 br_102 wl_47 vdd gnd cell_6t
Xbit_r48_c102 bl_102 br_102 wl_48 vdd gnd cell_6t
Xbit_r49_c102 bl_102 br_102 wl_49 vdd gnd cell_6t
Xbit_r50_c102 bl_102 br_102 wl_50 vdd gnd cell_6t
Xbit_r51_c102 bl_102 br_102 wl_51 vdd gnd cell_6t
Xbit_r52_c102 bl_102 br_102 wl_52 vdd gnd cell_6t
Xbit_r53_c102 bl_102 br_102 wl_53 vdd gnd cell_6t
Xbit_r54_c102 bl_102 br_102 wl_54 vdd gnd cell_6t
Xbit_r55_c102 bl_102 br_102 wl_55 vdd gnd cell_6t
Xbit_r56_c102 bl_102 br_102 wl_56 vdd gnd cell_6t
Xbit_r57_c102 bl_102 br_102 wl_57 vdd gnd cell_6t
Xbit_r58_c102 bl_102 br_102 wl_58 vdd gnd cell_6t
Xbit_r59_c102 bl_102 br_102 wl_59 vdd gnd cell_6t
Xbit_r60_c102 bl_102 br_102 wl_60 vdd gnd cell_6t
Xbit_r61_c102 bl_102 br_102 wl_61 vdd gnd cell_6t
Xbit_r62_c102 bl_102 br_102 wl_62 vdd gnd cell_6t
Xbit_r63_c102 bl_102 br_102 wl_63 vdd gnd cell_6t
Xbit_r64_c102 bl_102 br_102 wl_64 vdd gnd cell_6t
Xbit_r65_c102 bl_102 br_102 wl_65 vdd gnd cell_6t
Xbit_r66_c102 bl_102 br_102 wl_66 vdd gnd cell_6t
Xbit_r67_c102 bl_102 br_102 wl_67 vdd gnd cell_6t
Xbit_r68_c102 bl_102 br_102 wl_68 vdd gnd cell_6t
Xbit_r69_c102 bl_102 br_102 wl_69 vdd gnd cell_6t
Xbit_r70_c102 bl_102 br_102 wl_70 vdd gnd cell_6t
Xbit_r71_c102 bl_102 br_102 wl_71 vdd gnd cell_6t
Xbit_r72_c102 bl_102 br_102 wl_72 vdd gnd cell_6t
Xbit_r73_c102 bl_102 br_102 wl_73 vdd gnd cell_6t
Xbit_r74_c102 bl_102 br_102 wl_74 vdd gnd cell_6t
Xbit_r75_c102 bl_102 br_102 wl_75 vdd gnd cell_6t
Xbit_r76_c102 bl_102 br_102 wl_76 vdd gnd cell_6t
Xbit_r77_c102 bl_102 br_102 wl_77 vdd gnd cell_6t
Xbit_r78_c102 bl_102 br_102 wl_78 vdd gnd cell_6t
Xbit_r79_c102 bl_102 br_102 wl_79 vdd gnd cell_6t
Xbit_r80_c102 bl_102 br_102 wl_80 vdd gnd cell_6t
Xbit_r81_c102 bl_102 br_102 wl_81 vdd gnd cell_6t
Xbit_r82_c102 bl_102 br_102 wl_82 vdd gnd cell_6t
Xbit_r83_c102 bl_102 br_102 wl_83 vdd gnd cell_6t
Xbit_r84_c102 bl_102 br_102 wl_84 vdd gnd cell_6t
Xbit_r85_c102 bl_102 br_102 wl_85 vdd gnd cell_6t
Xbit_r86_c102 bl_102 br_102 wl_86 vdd gnd cell_6t
Xbit_r87_c102 bl_102 br_102 wl_87 vdd gnd cell_6t
Xbit_r88_c102 bl_102 br_102 wl_88 vdd gnd cell_6t
Xbit_r89_c102 bl_102 br_102 wl_89 vdd gnd cell_6t
Xbit_r90_c102 bl_102 br_102 wl_90 vdd gnd cell_6t
Xbit_r91_c102 bl_102 br_102 wl_91 vdd gnd cell_6t
Xbit_r92_c102 bl_102 br_102 wl_92 vdd gnd cell_6t
Xbit_r93_c102 bl_102 br_102 wl_93 vdd gnd cell_6t
Xbit_r94_c102 bl_102 br_102 wl_94 vdd gnd cell_6t
Xbit_r95_c102 bl_102 br_102 wl_95 vdd gnd cell_6t
Xbit_r96_c102 bl_102 br_102 wl_96 vdd gnd cell_6t
Xbit_r97_c102 bl_102 br_102 wl_97 vdd gnd cell_6t
Xbit_r98_c102 bl_102 br_102 wl_98 vdd gnd cell_6t
Xbit_r99_c102 bl_102 br_102 wl_99 vdd gnd cell_6t
Xbit_r100_c102 bl_102 br_102 wl_100 vdd gnd cell_6t
Xbit_r101_c102 bl_102 br_102 wl_101 vdd gnd cell_6t
Xbit_r102_c102 bl_102 br_102 wl_102 vdd gnd cell_6t
Xbit_r103_c102 bl_102 br_102 wl_103 vdd gnd cell_6t
Xbit_r104_c102 bl_102 br_102 wl_104 vdd gnd cell_6t
Xbit_r105_c102 bl_102 br_102 wl_105 vdd gnd cell_6t
Xbit_r106_c102 bl_102 br_102 wl_106 vdd gnd cell_6t
Xbit_r107_c102 bl_102 br_102 wl_107 vdd gnd cell_6t
Xbit_r108_c102 bl_102 br_102 wl_108 vdd gnd cell_6t
Xbit_r109_c102 bl_102 br_102 wl_109 vdd gnd cell_6t
Xbit_r110_c102 bl_102 br_102 wl_110 vdd gnd cell_6t
Xbit_r111_c102 bl_102 br_102 wl_111 vdd gnd cell_6t
Xbit_r112_c102 bl_102 br_102 wl_112 vdd gnd cell_6t
Xbit_r113_c102 bl_102 br_102 wl_113 vdd gnd cell_6t
Xbit_r114_c102 bl_102 br_102 wl_114 vdd gnd cell_6t
Xbit_r115_c102 bl_102 br_102 wl_115 vdd gnd cell_6t
Xbit_r116_c102 bl_102 br_102 wl_116 vdd gnd cell_6t
Xbit_r117_c102 bl_102 br_102 wl_117 vdd gnd cell_6t
Xbit_r118_c102 bl_102 br_102 wl_118 vdd gnd cell_6t
Xbit_r119_c102 bl_102 br_102 wl_119 vdd gnd cell_6t
Xbit_r120_c102 bl_102 br_102 wl_120 vdd gnd cell_6t
Xbit_r121_c102 bl_102 br_102 wl_121 vdd gnd cell_6t
Xbit_r122_c102 bl_102 br_102 wl_122 vdd gnd cell_6t
Xbit_r123_c102 bl_102 br_102 wl_123 vdd gnd cell_6t
Xbit_r124_c102 bl_102 br_102 wl_124 vdd gnd cell_6t
Xbit_r125_c102 bl_102 br_102 wl_125 vdd gnd cell_6t
Xbit_r126_c102 bl_102 br_102 wl_126 vdd gnd cell_6t
Xbit_r127_c102 bl_102 br_102 wl_127 vdd gnd cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd cell_6t
Xbit_r1_c103 bl_103 br_103 wl_1 vdd gnd cell_6t
Xbit_r2_c103 bl_103 br_103 wl_2 vdd gnd cell_6t
Xbit_r3_c103 bl_103 br_103 wl_3 vdd gnd cell_6t
Xbit_r4_c103 bl_103 br_103 wl_4 vdd gnd cell_6t
Xbit_r5_c103 bl_103 br_103 wl_5 vdd gnd cell_6t
Xbit_r6_c103 bl_103 br_103 wl_6 vdd gnd cell_6t
Xbit_r7_c103 bl_103 br_103 wl_7 vdd gnd cell_6t
Xbit_r8_c103 bl_103 br_103 wl_8 vdd gnd cell_6t
Xbit_r9_c103 bl_103 br_103 wl_9 vdd gnd cell_6t
Xbit_r10_c103 bl_103 br_103 wl_10 vdd gnd cell_6t
Xbit_r11_c103 bl_103 br_103 wl_11 vdd gnd cell_6t
Xbit_r12_c103 bl_103 br_103 wl_12 vdd gnd cell_6t
Xbit_r13_c103 bl_103 br_103 wl_13 vdd gnd cell_6t
Xbit_r14_c103 bl_103 br_103 wl_14 vdd gnd cell_6t
Xbit_r15_c103 bl_103 br_103 wl_15 vdd gnd cell_6t
Xbit_r16_c103 bl_103 br_103 wl_16 vdd gnd cell_6t
Xbit_r17_c103 bl_103 br_103 wl_17 vdd gnd cell_6t
Xbit_r18_c103 bl_103 br_103 wl_18 vdd gnd cell_6t
Xbit_r19_c103 bl_103 br_103 wl_19 vdd gnd cell_6t
Xbit_r20_c103 bl_103 br_103 wl_20 vdd gnd cell_6t
Xbit_r21_c103 bl_103 br_103 wl_21 vdd gnd cell_6t
Xbit_r22_c103 bl_103 br_103 wl_22 vdd gnd cell_6t
Xbit_r23_c103 bl_103 br_103 wl_23 vdd gnd cell_6t
Xbit_r24_c103 bl_103 br_103 wl_24 vdd gnd cell_6t
Xbit_r25_c103 bl_103 br_103 wl_25 vdd gnd cell_6t
Xbit_r26_c103 bl_103 br_103 wl_26 vdd gnd cell_6t
Xbit_r27_c103 bl_103 br_103 wl_27 vdd gnd cell_6t
Xbit_r28_c103 bl_103 br_103 wl_28 vdd gnd cell_6t
Xbit_r29_c103 bl_103 br_103 wl_29 vdd gnd cell_6t
Xbit_r30_c103 bl_103 br_103 wl_30 vdd gnd cell_6t
Xbit_r31_c103 bl_103 br_103 wl_31 vdd gnd cell_6t
Xbit_r32_c103 bl_103 br_103 wl_32 vdd gnd cell_6t
Xbit_r33_c103 bl_103 br_103 wl_33 vdd gnd cell_6t
Xbit_r34_c103 bl_103 br_103 wl_34 vdd gnd cell_6t
Xbit_r35_c103 bl_103 br_103 wl_35 vdd gnd cell_6t
Xbit_r36_c103 bl_103 br_103 wl_36 vdd gnd cell_6t
Xbit_r37_c103 bl_103 br_103 wl_37 vdd gnd cell_6t
Xbit_r38_c103 bl_103 br_103 wl_38 vdd gnd cell_6t
Xbit_r39_c103 bl_103 br_103 wl_39 vdd gnd cell_6t
Xbit_r40_c103 bl_103 br_103 wl_40 vdd gnd cell_6t
Xbit_r41_c103 bl_103 br_103 wl_41 vdd gnd cell_6t
Xbit_r42_c103 bl_103 br_103 wl_42 vdd gnd cell_6t
Xbit_r43_c103 bl_103 br_103 wl_43 vdd gnd cell_6t
Xbit_r44_c103 bl_103 br_103 wl_44 vdd gnd cell_6t
Xbit_r45_c103 bl_103 br_103 wl_45 vdd gnd cell_6t
Xbit_r46_c103 bl_103 br_103 wl_46 vdd gnd cell_6t
Xbit_r47_c103 bl_103 br_103 wl_47 vdd gnd cell_6t
Xbit_r48_c103 bl_103 br_103 wl_48 vdd gnd cell_6t
Xbit_r49_c103 bl_103 br_103 wl_49 vdd gnd cell_6t
Xbit_r50_c103 bl_103 br_103 wl_50 vdd gnd cell_6t
Xbit_r51_c103 bl_103 br_103 wl_51 vdd gnd cell_6t
Xbit_r52_c103 bl_103 br_103 wl_52 vdd gnd cell_6t
Xbit_r53_c103 bl_103 br_103 wl_53 vdd gnd cell_6t
Xbit_r54_c103 bl_103 br_103 wl_54 vdd gnd cell_6t
Xbit_r55_c103 bl_103 br_103 wl_55 vdd gnd cell_6t
Xbit_r56_c103 bl_103 br_103 wl_56 vdd gnd cell_6t
Xbit_r57_c103 bl_103 br_103 wl_57 vdd gnd cell_6t
Xbit_r58_c103 bl_103 br_103 wl_58 vdd gnd cell_6t
Xbit_r59_c103 bl_103 br_103 wl_59 vdd gnd cell_6t
Xbit_r60_c103 bl_103 br_103 wl_60 vdd gnd cell_6t
Xbit_r61_c103 bl_103 br_103 wl_61 vdd gnd cell_6t
Xbit_r62_c103 bl_103 br_103 wl_62 vdd gnd cell_6t
Xbit_r63_c103 bl_103 br_103 wl_63 vdd gnd cell_6t
Xbit_r64_c103 bl_103 br_103 wl_64 vdd gnd cell_6t
Xbit_r65_c103 bl_103 br_103 wl_65 vdd gnd cell_6t
Xbit_r66_c103 bl_103 br_103 wl_66 vdd gnd cell_6t
Xbit_r67_c103 bl_103 br_103 wl_67 vdd gnd cell_6t
Xbit_r68_c103 bl_103 br_103 wl_68 vdd gnd cell_6t
Xbit_r69_c103 bl_103 br_103 wl_69 vdd gnd cell_6t
Xbit_r70_c103 bl_103 br_103 wl_70 vdd gnd cell_6t
Xbit_r71_c103 bl_103 br_103 wl_71 vdd gnd cell_6t
Xbit_r72_c103 bl_103 br_103 wl_72 vdd gnd cell_6t
Xbit_r73_c103 bl_103 br_103 wl_73 vdd gnd cell_6t
Xbit_r74_c103 bl_103 br_103 wl_74 vdd gnd cell_6t
Xbit_r75_c103 bl_103 br_103 wl_75 vdd gnd cell_6t
Xbit_r76_c103 bl_103 br_103 wl_76 vdd gnd cell_6t
Xbit_r77_c103 bl_103 br_103 wl_77 vdd gnd cell_6t
Xbit_r78_c103 bl_103 br_103 wl_78 vdd gnd cell_6t
Xbit_r79_c103 bl_103 br_103 wl_79 vdd gnd cell_6t
Xbit_r80_c103 bl_103 br_103 wl_80 vdd gnd cell_6t
Xbit_r81_c103 bl_103 br_103 wl_81 vdd gnd cell_6t
Xbit_r82_c103 bl_103 br_103 wl_82 vdd gnd cell_6t
Xbit_r83_c103 bl_103 br_103 wl_83 vdd gnd cell_6t
Xbit_r84_c103 bl_103 br_103 wl_84 vdd gnd cell_6t
Xbit_r85_c103 bl_103 br_103 wl_85 vdd gnd cell_6t
Xbit_r86_c103 bl_103 br_103 wl_86 vdd gnd cell_6t
Xbit_r87_c103 bl_103 br_103 wl_87 vdd gnd cell_6t
Xbit_r88_c103 bl_103 br_103 wl_88 vdd gnd cell_6t
Xbit_r89_c103 bl_103 br_103 wl_89 vdd gnd cell_6t
Xbit_r90_c103 bl_103 br_103 wl_90 vdd gnd cell_6t
Xbit_r91_c103 bl_103 br_103 wl_91 vdd gnd cell_6t
Xbit_r92_c103 bl_103 br_103 wl_92 vdd gnd cell_6t
Xbit_r93_c103 bl_103 br_103 wl_93 vdd gnd cell_6t
Xbit_r94_c103 bl_103 br_103 wl_94 vdd gnd cell_6t
Xbit_r95_c103 bl_103 br_103 wl_95 vdd gnd cell_6t
Xbit_r96_c103 bl_103 br_103 wl_96 vdd gnd cell_6t
Xbit_r97_c103 bl_103 br_103 wl_97 vdd gnd cell_6t
Xbit_r98_c103 bl_103 br_103 wl_98 vdd gnd cell_6t
Xbit_r99_c103 bl_103 br_103 wl_99 vdd gnd cell_6t
Xbit_r100_c103 bl_103 br_103 wl_100 vdd gnd cell_6t
Xbit_r101_c103 bl_103 br_103 wl_101 vdd gnd cell_6t
Xbit_r102_c103 bl_103 br_103 wl_102 vdd gnd cell_6t
Xbit_r103_c103 bl_103 br_103 wl_103 vdd gnd cell_6t
Xbit_r104_c103 bl_103 br_103 wl_104 vdd gnd cell_6t
Xbit_r105_c103 bl_103 br_103 wl_105 vdd gnd cell_6t
Xbit_r106_c103 bl_103 br_103 wl_106 vdd gnd cell_6t
Xbit_r107_c103 bl_103 br_103 wl_107 vdd gnd cell_6t
Xbit_r108_c103 bl_103 br_103 wl_108 vdd gnd cell_6t
Xbit_r109_c103 bl_103 br_103 wl_109 vdd gnd cell_6t
Xbit_r110_c103 bl_103 br_103 wl_110 vdd gnd cell_6t
Xbit_r111_c103 bl_103 br_103 wl_111 vdd gnd cell_6t
Xbit_r112_c103 bl_103 br_103 wl_112 vdd gnd cell_6t
Xbit_r113_c103 bl_103 br_103 wl_113 vdd gnd cell_6t
Xbit_r114_c103 bl_103 br_103 wl_114 vdd gnd cell_6t
Xbit_r115_c103 bl_103 br_103 wl_115 vdd gnd cell_6t
Xbit_r116_c103 bl_103 br_103 wl_116 vdd gnd cell_6t
Xbit_r117_c103 bl_103 br_103 wl_117 vdd gnd cell_6t
Xbit_r118_c103 bl_103 br_103 wl_118 vdd gnd cell_6t
Xbit_r119_c103 bl_103 br_103 wl_119 vdd gnd cell_6t
Xbit_r120_c103 bl_103 br_103 wl_120 vdd gnd cell_6t
Xbit_r121_c103 bl_103 br_103 wl_121 vdd gnd cell_6t
Xbit_r122_c103 bl_103 br_103 wl_122 vdd gnd cell_6t
Xbit_r123_c103 bl_103 br_103 wl_123 vdd gnd cell_6t
Xbit_r124_c103 bl_103 br_103 wl_124 vdd gnd cell_6t
Xbit_r125_c103 bl_103 br_103 wl_125 vdd gnd cell_6t
Xbit_r126_c103 bl_103 br_103 wl_126 vdd gnd cell_6t
Xbit_r127_c103 bl_103 br_103 wl_127 vdd gnd cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd cell_6t
Xbit_r1_c104 bl_104 br_104 wl_1 vdd gnd cell_6t
Xbit_r2_c104 bl_104 br_104 wl_2 vdd gnd cell_6t
Xbit_r3_c104 bl_104 br_104 wl_3 vdd gnd cell_6t
Xbit_r4_c104 bl_104 br_104 wl_4 vdd gnd cell_6t
Xbit_r5_c104 bl_104 br_104 wl_5 vdd gnd cell_6t
Xbit_r6_c104 bl_104 br_104 wl_6 vdd gnd cell_6t
Xbit_r7_c104 bl_104 br_104 wl_7 vdd gnd cell_6t
Xbit_r8_c104 bl_104 br_104 wl_8 vdd gnd cell_6t
Xbit_r9_c104 bl_104 br_104 wl_9 vdd gnd cell_6t
Xbit_r10_c104 bl_104 br_104 wl_10 vdd gnd cell_6t
Xbit_r11_c104 bl_104 br_104 wl_11 vdd gnd cell_6t
Xbit_r12_c104 bl_104 br_104 wl_12 vdd gnd cell_6t
Xbit_r13_c104 bl_104 br_104 wl_13 vdd gnd cell_6t
Xbit_r14_c104 bl_104 br_104 wl_14 vdd gnd cell_6t
Xbit_r15_c104 bl_104 br_104 wl_15 vdd gnd cell_6t
Xbit_r16_c104 bl_104 br_104 wl_16 vdd gnd cell_6t
Xbit_r17_c104 bl_104 br_104 wl_17 vdd gnd cell_6t
Xbit_r18_c104 bl_104 br_104 wl_18 vdd gnd cell_6t
Xbit_r19_c104 bl_104 br_104 wl_19 vdd gnd cell_6t
Xbit_r20_c104 bl_104 br_104 wl_20 vdd gnd cell_6t
Xbit_r21_c104 bl_104 br_104 wl_21 vdd gnd cell_6t
Xbit_r22_c104 bl_104 br_104 wl_22 vdd gnd cell_6t
Xbit_r23_c104 bl_104 br_104 wl_23 vdd gnd cell_6t
Xbit_r24_c104 bl_104 br_104 wl_24 vdd gnd cell_6t
Xbit_r25_c104 bl_104 br_104 wl_25 vdd gnd cell_6t
Xbit_r26_c104 bl_104 br_104 wl_26 vdd gnd cell_6t
Xbit_r27_c104 bl_104 br_104 wl_27 vdd gnd cell_6t
Xbit_r28_c104 bl_104 br_104 wl_28 vdd gnd cell_6t
Xbit_r29_c104 bl_104 br_104 wl_29 vdd gnd cell_6t
Xbit_r30_c104 bl_104 br_104 wl_30 vdd gnd cell_6t
Xbit_r31_c104 bl_104 br_104 wl_31 vdd gnd cell_6t
Xbit_r32_c104 bl_104 br_104 wl_32 vdd gnd cell_6t
Xbit_r33_c104 bl_104 br_104 wl_33 vdd gnd cell_6t
Xbit_r34_c104 bl_104 br_104 wl_34 vdd gnd cell_6t
Xbit_r35_c104 bl_104 br_104 wl_35 vdd gnd cell_6t
Xbit_r36_c104 bl_104 br_104 wl_36 vdd gnd cell_6t
Xbit_r37_c104 bl_104 br_104 wl_37 vdd gnd cell_6t
Xbit_r38_c104 bl_104 br_104 wl_38 vdd gnd cell_6t
Xbit_r39_c104 bl_104 br_104 wl_39 vdd gnd cell_6t
Xbit_r40_c104 bl_104 br_104 wl_40 vdd gnd cell_6t
Xbit_r41_c104 bl_104 br_104 wl_41 vdd gnd cell_6t
Xbit_r42_c104 bl_104 br_104 wl_42 vdd gnd cell_6t
Xbit_r43_c104 bl_104 br_104 wl_43 vdd gnd cell_6t
Xbit_r44_c104 bl_104 br_104 wl_44 vdd gnd cell_6t
Xbit_r45_c104 bl_104 br_104 wl_45 vdd gnd cell_6t
Xbit_r46_c104 bl_104 br_104 wl_46 vdd gnd cell_6t
Xbit_r47_c104 bl_104 br_104 wl_47 vdd gnd cell_6t
Xbit_r48_c104 bl_104 br_104 wl_48 vdd gnd cell_6t
Xbit_r49_c104 bl_104 br_104 wl_49 vdd gnd cell_6t
Xbit_r50_c104 bl_104 br_104 wl_50 vdd gnd cell_6t
Xbit_r51_c104 bl_104 br_104 wl_51 vdd gnd cell_6t
Xbit_r52_c104 bl_104 br_104 wl_52 vdd gnd cell_6t
Xbit_r53_c104 bl_104 br_104 wl_53 vdd gnd cell_6t
Xbit_r54_c104 bl_104 br_104 wl_54 vdd gnd cell_6t
Xbit_r55_c104 bl_104 br_104 wl_55 vdd gnd cell_6t
Xbit_r56_c104 bl_104 br_104 wl_56 vdd gnd cell_6t
Xbit_r57_c104 bl_104 br_104 wl_57 vdd gnd cell_6t
Xbit_r58_c104 bl_104 br_104 wl_58 vdd gnd cell_6t
Xbit_r59_c104 bl_104 br_104 wl_59 vdd gnd cell_6t
Xbit_r60_c104 bl_104 br_104 wl_60 vdd gnd cell_6t
Xbit_r61_c104 bl_104 br_104 wl_61 vdd gnd cell_6t
Xbit_r62_c104 bl_104 br_104 wl_62 vdd gnd cell_6t
Xbit_r63_c104 bl_104 br_104 wl_63 vdd gnd cell_6t
Xbit_r64_c104 bl_104 br_104 wl_64 vdd gnd cell_6t
Xbit_r65_c104 bl_104 br_104 wl_65 vdd gnd cell_6t
Xbit_r66_c104 bl_104 br_104 wl_66 vdd gnd cell_6t
Xbit_r67_c104 bl_104 br_104 wl_67 vdd gnd cell_6t
Xbit_r68_c104 bl_104 br_104 wl_68 vdd gnd cell_6t
Xbit_r69_c104 bl_104 br_104 wl_69 vdd gnd cell_6t
Xbit_r70_c104 bl_104 br_104 wl_70 vdd gnd cell_6t
Xbit_r71_c104 bl_104 br_104 wl_71 vdd gnd cell_6t
Xbit_r72_c104 bl_104 br_104 wl_72 vdd gnd cell_6t
Xbit_r73_c104 bl_104 br_104 wl_73 vdd gnd cell_6t
Xbit_r74_c104 bl_104 br_104 wl_74 vdd gnd cell_6t
Xbit_r75_c104 bl_104 br_104 wl_75 vdd gnd cell_6t
Xbit_r76_c104 bl_104 br_104 wl_76 vdd gnd cell_6t
Xbit_r77_c104 bl_104 br_104 wl_77 vdd gnd cell_6t
Xbit_r78_c104 bl_104 br_104 wl_78 vdd gnd cell_6t
Xbit_r79_c104 bl_104 br_104 wl_79 vdd gnd cell_6t
Xbit_r80_c104 bl_104 br_104 wl_80 vdd gnd cell_6t
Xbit_r81_c104 bl_104 br_104 wl_81 vdd gnd cell_6t
Xbit_r82_c104 bl_104 br_104 wl_82 vdd gnd cell_6t
Xbit_r83_c104 bl_104 br_104 wl_83 vdd gnd cell_6t
Xbit_r84_c104 bl_104 br_104 wl_84 vdd gnd cell_6t
Xbit_r85_c104 bl_104 br_104 wl_85 vdd gnd cell_6t
Xbit_r86_c104 bl_104 br_104 wl_86 vdd gnd cell_6t
Xbit_r87_c104 bl_104 br_104 wl_87 vdd gnd cell_6t
Xbit_r88_c104 bl_104 br_104 wl_88 vdd gnd cell_6t
Xbit_r89_c104 bl_104 br_104 wl_89 vdd gnd cell_6t
Xbit_r90_c104 bl_104 br_104 wl_90 vdd gnd cell_6t
Xbit_r91_c104 bl_104 br_104 wl_91 vdd gnd cell_6t
Xbit_r92_c104 bl_104 br_104 wl_92 vdd gnd cell_6t
Xbit_r93_c104 bl_104 br_104 wl_93 vdd gnd cell_6t
Xbit_r94_c104 bl_104 br_104 wl_94 vdd gnd cell_6t
Xbit_r95_c104 bl_104 br_104 wl_95 vdd gnd cell_6t
Xbit_r96_c104 bl_104 br_104 wl_96 vdd gnd cell_6t
Xbit_r97_c104 bl_104 br_104 wl_97 vdd gnd cell_6t
Xbit_r98_c104 bl_104 br_104 wl_98 vdd gnd cell_6t
Xbit_r99_c104 bl_104 br_104 wl_99 vdd gnd cell_6t
Xbit_r100_c104 bl_104 br_104 wl_100 vdd gnd cell_6t
Xbit_r101_c104 bl_104 br_104 wl_101 vdd gnd cell_6t
Xbit_r102_c104 bl_104 br_104 wl_102 vdd gnd cell_6t
Xbit_r103_c104 bl_104 br_104 wl_103 vdd gnd cell_6t
Xbit_r104_c104 bl_104 br_104 wl_104 vdd gnd cell_6t
Xbit_r105_c104 bl_104 br_104 wl_105 vdd gnd cell_6t
Xbit_r106_c104 bl_104 br_104 wl_106 vdd gnd cell_6t
Xbit_r107_c104 bl_104 br_104 wl_107 vdd gnd cell_6t
Xbit_r108_c104 bl_104 br_104 wl_108 vdd gnd cell_6t
Xbit_r109_c104 bl_104 br_104 wl_109 vdd gnd cell_6t
Xbit_r110_c104 bl_104 br_104 wl_110 vdd gnd cell_6t
Xbit_r111_c104 bl_104 br_104 wl_111 vdd gnd cell_6t
Xbit_r112_c104 bl_104 br_104 wl_112 vdd gnd cell_6t
Xbit_r113_c104 bl_104 br_104 wl_113 vdd gnd cell_6t
Xbit_r114_c104 bl_104 br_104 wl_114 vdd gnd cell_6t
Xbit_r115_c104 bl_104 br_104 wl_115 vdd gnd cell_6t
Xbit_r116_c104 bl_104 br_104 wl_116 vdd gnd cell_6t
Xbit_r117_c104 bl_104 br_104 wl_117 vdd gnd cell_6t
Xbit_r118_c104 bl_104 br_104 wl_118 vdd gnd cell_6t
Xbit_r119_c104 bl_104 br_104 wl_119 vdd gnd cell_6t
Xbit_r120_c104 bl_104 br_104 wl_120 vdd gnd cell_6t
Xbit_r121_c104 bl_104 br_104 wl_121 vdd gnd cell_6t
Xbit_r122_c104 bl_104 br_104 wl_122 vdd gnd cell_6t
Xbit_r123_c104 bl_104 br_104 wl_123 vdd gnd cell_6t
Xbit_r124_c104 bl_104 br_104 wl_124 vdd gnd cell_6t
Xbit_r125_c104 bl_104 br_104 wl_125 vdd gnd cell_6t
Xbit_r126_c104 bl_104 br_104 wl_126 vdd gnd cell_6t
Xbit_r127_c104 bl_104 br_104 wl_127 vdd gnd cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd cell_6t
Xbit_r1_c105 bl_105 br_105 wl_1 vdd gnd cell_6t
Xbit_r2_c105 bl_105 br_105 wl_2 vdd gnd cell_6t
Xbit_r3_c105 bl_105 br_105 wl_3 vdd gnd cell_6t
Xbit_r4_c105 bl_105 br_105 wl_4 vdd gnd cell_6t
Xbit_r5_c105 bl_105 br_105 wl_5 vdd gnd cell_6t
Xbit_r6_c105 bl_105 br_105 wl_6 vdd gnd cell_6t
Xbit_r7_c105 bl_105 br_105 wl_7 vdd gnd cell_6t
Xbit_r8_c105 bl_105 br_105 wl_8 vdd gnd cell_6t
Xbit_r9_c105 bl_105 br_105 wl_9 vdd gnd cell_6t
Xbit_r10_c105 bl_105 br_105 wl_10 vdd gnd cell_6t
Xbit_r11_c105 bl_105 br_105 wl_11 vdd gnd cell_6t
Xbit_r12_c105 bl_105 br_105 wl_12 vdd gnd cell_6t
Xbit_r13_c105 bl_105 br_105 wl_13 vdd gnd cell_6t
Xbit_r14_c105 bl_105 br_105 wl_14 vdd gnd cell_6t
Xbit_r15_c105 bl_105 br_105 wl_15 vdd gnd cell_6t
Xbit_r16_c105 bl_105 br_105 wl_16 vdd gnd cell_6t
Xbit_r17_c105 bl_105 br_105 wl_17 vdd gnd cell_6t
Xbit_r18_c105 bl_105 br_105 wl_18 vdd gnd cell_6t
Xbit_r19_c105 bl_105 br_105 wl_19 vdd gnd cell_6t
Xbit_r20_c105 bl_105 br_105 wl_20 vdd gnd cell_6t
Xbit_r21_c105 bl_105 br_105 wl_21 vdd gnd cell_6t
Xbit_r22_c105 bl_105 br_105 wl_22 vdd gnd cell_6t
Xbit_r23_c105 bl_105 br_105 wl_23 vdd gnd cell_6t
Xbit_r24_c105 bl_105 br_105 wl_24 vdd gnd cell_6t
Xbit_r25_c105 bl_105 br_105 wl_25 vdd gnd cell_6t
Xbit_r26_c105 bl_105 br_105 wl_26 vdd gnd cell_6t
Xbit_r27_c105 bl_105 br_105 wl_27 vdd gnd cell_6t
Xbit_r28_c105 bl_105 br_105 wl_28 vdd gnd cell_6t
Xbit_r29_c105 bl_105 br_105 wl_29 vdd gnd cell_6t
Xbit_r30_c105 bl_105 br_105 wl_30 vdd gnd cell_6t
Xbit_r31_c105 bl_105 br_105 wl_31 vdd gnd cell_6t
Xbit_r32_c105 bl_105 br_105 wl_32 vdd gnd cell_6t
Xbit_r33_c105 bl_105 br_105 wl_33 vdd gnd cell_6t
Xbit_r34_c105 bl_105 br_105 wl_34 vdd gnd cell_6t
Xbit_r35_c105 bl_105 br_105 wl_35 vdd gnd cell_6t
Xbit_r36_c105 bl_105 br_105 wl_36 vdd gnd cell_6t
Xbit_r37_c105 bl_105 br_105 wl_37 vdd gnd cell_6t
Xbit_r38_c105 bl_105 br_105 wl_38 vdd gnd cell_6t
Xbit_r39_c105 bl_105 br_105 wl_39 vdd gnd cell_6t
Xbit_r40_c105 bl_105 br_105 wl_40 vdd gnd cell_6t
Xbit_r41_c105 bl_105 br_105 wl_41 vdd gnd cell_6t
Xbit_r42_c105 bl_105 br_105 wl_42 vdd gnd cell_6t
Xbit_r43_c105 bl_105 br_105 wl_43 vdd gnd cell_6t
Xbit_r44_c105 bl_105 br_105 wl_44 vdd gnd cell_6t
Xbit_r45_c105 bl_105 br_105 wl_45 vdd gnd cell_6t
Xbit_r46_c105 bl_105 br_105 wl_46 vdd gnd cell_6t
Xbit_r47_c105 bl_105 br_105 wl_47 vdd gnd cell_6t
Xbit_r48_c105 bl_105 br_105 wl_48 vdd gnd cell_6t
Xbit_r49_c105 bl_105 br_105 wl_49 vdd gnd cell_6t
Xbit_r50_c105 bl_105 br_105 wl_50 vdd gnd cell_6t
Xbit_r51_c105 bl_105 br_105 wl_51 vdd gnd cell_6t
Xbit_r52_c105 bl_105 br_105 wl_52 vdd gnd cell_6t
Xbit_r53_c105 bl_105 br_105 wl_53 vdd gnd cell_6t
Xbit_r54_c105 bl_105 br_105 wl_54 vdd gnd cell_6t
Xbit_r55_c105 bl_105 br_105 wl_55 vdd gnd cell_6t
Xbit_r56_c105 bl_105 br_105 wl_56 vdd gnd cell_6t
Xbit_r57_c105 bl_105 br_105 wl_57 vdd gnd cell_6t
Xbit_r58_c105 bl_105 br_105 wl_58 vdd gnd cell_6t
Xbit_r59_c105 bl_105 br_105 wl_59 vdd gnd cell_6t
Xbit_r60_c105 bl_105 br_105 wl_60 vdd gnd cell_6t
Xbit_r61_c105 bl_105 br_105 wl_61 vdd gnd cell_6t
Xbit_r62_c105 bl_105 br_105 wl_62 vdd gnd cell_6t
Xbit_r63_c105 bl_105 br_105 wl_63 vdd gnd cell_6t
Xbit_r64_c105 bl_105 br_105 wl_64 vdd gnd cell_6t
Xbit_r65_c105 bl_105 br_105 wl_65 vdd gnd cell_6t
Xbit_r66_c105 bl_105 br_105 wl_66 vdd gnd cell_6t
Xbit_r67_c105 bl_105 br_105 wl_67 vdd gnd cell_6t
Xbit_r68_c105 bl_105 br_105 wl_68 vdd gnd cell_6t
Xbit_r69_c105 bl_105 br_105 wl_69 vdd gnd cell_6t
Xbit_r70_c105 bl_105 br_105 wl_70 vdd gnd cell_6t
Xbit_r71_c105 bl_105 br_105 wl_71 vdd gnd cell_6t
Xbit_r72_c105 bl_105 br_105 wl_72 vdd gnd cell_6t
Xbit_r73_c105 bl_105 br_105 wl_73 vdd gnd cell_6t
Xbit_r74_c105 bl_105 br_105 wl_74 vdd gnd cell_6t
Xbit_r75_c105 bl_105 br_105 wl_75 vdd gnd cell_6t
Xbit_r76_c105 bl_105 br_105 wl_76 vdd gnd cell_6t
Xbit_r77_c105 bl_105 br_105 wl_77 vdd gnd cell_6t
Xbit_r78_c105 bl_105 br_105 wl_78 vdd gnd cell_6t
Xbit_r79_c105 bl_105 br_105 wl_79 vdd gnd cell_6t
Xbit_r80_c105 bl_105 br_105 wl_80 vdd gnd cell_6t
Xbit_r81_c105 bl_105 br_105 wl_81 vdd gnd cell_6t
Xbit_r82_c105 bl_105 br_105 wl_82 vdd gnd cell_6t
Xbit_r83_c105 bl_105 br_105 wl_83 vdd gnd cell_6t
Xbit_r84_c105 bl_105 br_105 wl_84 vdd gnd cell_6t
Xbit_r85_c105 bl_105 br_105 wl_85 vdd gnd cell_6t
Xbit_r86_c105 bl_105 br_105 wl_86 vdd gnd cell_6t
Xbit_r87_c105 bl_105 br_105 wl_87 vdd gnd cell_6t
Xbit_r88_c105 bl_105 br_105 wl_88 vdd gnd cell_6t
Xbit_r89_c105 bl_105 br_105 wl_89 vdd gnd cell_6t
Xbit_r90_c105 bl_105 br_105 wl_90 vdd gnd cell_6t
Xbit_r91_c105 bl_105 br_105 wl_91 vdd gnd cell_6t
Xbit_r92_c105 bl_105 br_105 wl_92 vdd gnd cell_6t
Xbit_r93_c105 bl_105 br_105 wl_93 vdd gnd cell_6t
Xbit_r94_c105 bl_105 br_105 wl_94 vdd gnd cell_6t
Xbit_r95_c105 bl_105 br_105 wl_95 vdd gnd cell_6t
Xbit_r96_c105 bl_105 br_105 wl_96 vdd gnd cell_6t
Xbit_r97_c105 bl_105 br_105 wl_97 vdd gnd cell_6t
Xbit_r98_c105 bl_105 br_105 wl_98 vdd gnd cell_6t
Xbit_r99_c105 bl_105 br_105 wl_99 vdd gnd cell_6t
Xbit_r100_c105 bl_105 br_105 wl_100 vdd gnd cell_6t
Xbit_r101_c105 bl_105 br_105 wl_101 vdd gnd cell_6t
Xbit_r102_c105 bl_105 br_105 wl_102 vdd gnd cell_6t
Xbit_r103_c105 bl_105 br_105 wl_103 vdd gnd cell_6t
Xbit_r104_c105 bl_105 br_105 wl_104 vdd gnd cell_6t
Xbit_r105_c105 bl_105 br_105 wl_105 vdd gnd cell_6t
Xbit_r106_c105 bl_105 br_105 wl_106 vdd gnd cell_6t
Xbit_r107_c105 bl_105 br_105 wl_107 vdd gnd cell_6t
Xbit_r108_c105 bl_105 br_105 wl_108 vdd gnd cell_6t
Xbit_r109_c105 bl_105 br_105 wl_109 vdd gnd cell_6t
Xbit_r110_c105 bl_105 br_105 wl_110 vdd gnd cell_6t
Xbit_r111_c105 bl_105 br_105 wl_111 vdd gnd cell_6t
Xbit_r112_c105 bl_105 br_105 wl_112 vdd gnd cell_6t
Xbit_r113_c105 bl_105 br_105 wl_113 vdd gnd cell_6t
Xbit_r114_c105 bl_105 br_105 wl_114 vdd gnd cell_6t
Xbit_r115_c105 bl_105 br_105 wl_115 vdd gnd cell_6t
Xbit_r116_c105 bl_105 br_105 wl_116 vdd gnd cell_6t
Xbit_r117_c105 bl_105 br_105 wl_117 vdd gnd cell_6t
Xbit_r118_c105 bl_105 br_105 wl_118 vdd gnd cell_6t
Xbit_r119_c105 bl_105 br_105 wl_119 vdd gnd cell_6t
Xbit_r120_c105 bl_105 br_105 wl_120 vdd gnd cell_6t
Xbit_r121_c105 bl_105 br_105 wl_121 vdd gnd cell_6t
Xbit_r122_c105 bl_105 br_105 wl_122 vdd gnd cell_6t
Xbit_r123_c105 bl_105 br_105 wl_123 vdd gnd cell_6t
Xbit_r124_c105 bl_105 br_105 wl_124 vdd gnd cell_6t
Xbit_r125_c105 bl_105 br_105 wl_125 vdd gnd cell_6t
Xbit_r126_c105 bl_105 br_105 wl_126 vdd gnd cell_6t
Xbit_r127_c105 bl_105 br_105 wl_127 vdd gnd cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd cell_6t
Xbit_r1_c106 bl_106 br_106 wl_1 vdd gnd cell_6t
Xbit_r2_c106 bl_106 br_106 wl_2 vdd gnd cell_6t
Xbit_r3_c106 bl_106 br_106 wl_3 vdd gnd cell_6t
Xbit_r4_c106 bl_106 br_106 wl_4 vdd gnd cell_6t
Xbit_r5_c106 bl_106 br_106 wl_5 vdd gnd cell_6t
Xbit_r6_c106 bl_106 br_106 wl_6 vdd gnd cell_6t
Xbit_r7_c106 bl_106 br_106 wl_7 vdd gnd cell_6t
Xbit_r8_c106 bl_106 br_106 wl_8 vdd gnd cell_6t
Xbit_r9_c106 bl_106 br_106 wl_9 vdd gnd cell_6t
Xbit_r10_c106 bl_106 br_106 wl_10 vdd gnd cell_6t
Xbit_r11_c106 bl_106 br_106 wl_11 vdd gnd cell_6t
Xbit_r12_c106 bl_106 br_106 wl_12 vdd gnd cell_6t
Xbit_r13_c106 bl_106 br_106 wl_13 vdd gnd cell_6t
Xbit_r14_c106 bl_106 br_106 wl_14 vdd gnd cell_6t
Xbit_r15_c106 bl_106 br_106 wl_15 vdd gnd cell_6t
Xbit_r16_c106 bl_106 br_106 wl_16 vdd gnd cell_6t
Xbit_r17_c106 bl_106 br_106 wl_17 vdd gnd cell_6t
Xbit_r18_c106 bl_106 br_106 wl_18 vdd gnd cell_6t
Xbit_r19_c106 bl_106 br_106 wl_19 vdd gnd cell_6t
Xbit_r20_c106 bl_106 br_106 wl_20 vdd gnd cell_6t
Xbit_r21_c106 bl_106 br_106 wl_21 vdd gnd cell_6t
Xbit_r22_c106 bl_106 br_106 wl_22 vdd gnd cell_6t
Xbit_r23_c106 bl_106 br_106 wl_23 vdd gnd cell_6t
Xbit_r24_c106 bl_106 br_106 wl_24 vdd gnd cell_6t
Xbit_r25_c106 bl_106 br_106 wl_25 vdd gnd cell_6t
Xbit_r26_c106 bl_106 br_106 wl_26 vdd gnd cell_6t
Xbit_r27_c106 bl_106 br_106 wl_27 vdd gnd cell_6t
Xbit_r28_c106 bl_106 br_106 wl_28 vdd gnd cell_6t
Xbit_r29_c106 bl_106 br_106 wl_29 vdd gnd cell_6t
Xbit_r30_c106 bl_106 br_106 wl_30 vdd gnd cell_6t
Xbit_r31_c106 bl_106 br_106 wl_31 vdd gnd cell_6t
Xbit_r32_c106 bl_106 br_106 wl_32 vdd gnd cell_6t
Xbit_r33_c106 bl_106 br_106 wl_33 vdd gnd cell_6t
Xbit_r34_c106 bl_106 br_106 wl_34 vdd gnd cell_6t
Xbit_r35_c106 bl_106 br_106 wl_35 vdd gnd cell_6t
Xbit_r36_c106 bl_106 br_106 wl_36 vdd gnd cell_6t
Xbit_r37_c106 bl_106 br_106 wl_37 vdd gnd cell_6t
Xbit_r38_c106 bl_106 br_106 wl_38 vdd gnd cell_6t
Xbit_r39_c106 bl_106 br_106 wl_39 vdd gnd cell_6t
Xbit_r40_c106 bl_106 br_106 wl_40 vdd gnd cell_6t
Xbit_r41_c106 bl_106 br_106 wl_41 vdd gnd cell_6t
Xbit_r42_c106 bl_106 br_106 wl_42 vdd gnd cell_6t
Xbit_r43_c106 bl_106 br_106 wl_43 vdd gnd cell_6t
Xbit_r44_c106 bl_106 br_106 wl_44 vdd gnd cell_6t
Xbit_r45_c106 bl_106 br_106 wl_45 vdd gnd cell_6t
Xbit_r46_c106 bl_106 br_106 wl_46 vdd gnd cell_6t
Xbit_r47_c106 bl_106 br_106 wl_47 vdd gnd cell_6t
Xbit_r48_c106 bl_106 br_106 wl_48 vdd gnd cell_6t
Xbit_r49_c106 bl_106 br_106 wl_49 vdd gnd cell_6t
Xbit_r50_c106 bl_106 br_106 wl_50 vdd gnd cell_6t
Xbit_r51_c106 bl_106 br_106 wl_51 vdd gnd cell_6t
Xbit_r52_c106 bl_106 br_106 wl_52 vdd gnd cell_6t
Xbit_r53_c106 bl_106 br_106 wl_53 vdd gnd cell_6t
Xbit_r54_c106 bl_106 br_106 wl_54 vdd gnd cell_6t
Xbit_r55_c106 bl_106 br_106 wl_55 vdd gnd cell_6t
Xbit_r56_c106 bl_106 br_106 wl_56 vdd gnd cell_6t
Xbit_r57_c106 bl_106 br_106 wl_57 vdd gnd cell_6t
Xbit_r58_c106 bl_106 br_106 wl_58 vdd gnd cell_6t
Xbit_r59_c106 bl_106 br_106 wl_59 vdd gnd cell_6t
Xbit_r60_c106 bl_106 br_106 wl_60 vdd gnd cell_6t
Xbit_r61_c106 bl_106 br_106 wl_61 vdd gnd cell_6t
Xbit_r62_c106 bl_106 br_106 wl_62 vdd gnd cell_6t
Xbit_r63_c106 bl_106 br_106 wl_63 vdd gnd cell_6t
Xbit_r64_c106 bl_106 br_106 wl_64 vdd gnd cell_6t
Xbit_r65_c106 bl_106 br_106 wl_65 vdd gnd cell_6t
Xbit_r66_c106 bl_106 br_106 wl_66 vdd gnd cell_6t
Xbit_r67_c106 bl_106 br_106 wl_67 vdd gnd cell_6t
Xbit_r68_c106 bl_106 br_106 wl_68 vdd gnd cell_6t
Xbit_r69_c106 bl_106 br_106 wl_69 vdd gnd cell_6t
Xbit_r70_c106 bl_106 br_106 wl_70 vdd gnd cell_6t
Xbit_r71_c106 bl_106 br_106 wl_71 vdd gnd cell_6t
Xbit_r72_c106 bl_106 br_106 wl_72 vdd gnd cell_6t
Xbit_r73_c106 bl_106 br_106 wl_73 vdd gnd cell_6t
Xbit_r74_c106 bl_106 br_106 wl_74 vdd gnd cell_6t
Xbit_r75_c106 bl_106 br_106 wl_75 vdd gnd cell_6t
Xbit_r76_c106 bl_106 br_106 wl_76 vdd gnd cell_6t
Xbit_r77_c106 bl_106 br_106 wl_77 vdd gnd cell_6t
Xbit_r78_c106 bl_106 br_106 wl_78 vdd gnd cell_6t
Xbit_r79_c106 bl_106 br_106 wl_79 vdd gnd cell_6t
Xbit_r80_c106 bl_106 br_106 wl_80 vdd gnd cell_6t
Xbit_r81_c106 bl_106 br_106 wl_81 vdd gnd cell_6t
Xbit_r82_c106 bl_106 br_106 wl_82 vdd gnd cell_6t
Xbit_r83_c106 bl_106 br_106 wl_83 vdd gnd cell_6t
Xbit_r84_c106 bl_106 br_106 wl_84 vdd gnd cell_6t
Xbit_r85_c106 bl_106 br_106 wl_85 vdd gnd cell_6t
Xbit_r86_c106 bl_106 br_106 wl_86 vdd gnd cell_6t
Xbit_r87_c106 bl_106 br_106 wl_87 vdd gnd cell_6t
Xbit_r88_c106 bl_106 br_106 wl_88 vdd gnd cell_6t
Xbit_r89_c106 bl_106 br_106 wl_89 vdd gnd cell_6t
Xbit_r90_c106 bl_106 br_106 wl_90 vdd gnd cell_6t
Xbit_r91_c106 bl_106 br_106 wl_91 vdd gnd cell_6t
Xbit_r92_c106 bl_106 br_106 wl_92 vdd gnd cell_6t
Xbit_r93_c106 bl_106 br_106 wl_93 vdd gnd cell_6t
Xbit_r94_c106 bl_106 br_106 wl_94 vdd gnd cell_6t
Xbit_r95_c106 bl_106 br_106 wl_95 vdd gnd cell_6t
Xbit_r96_c106 bl_106 br_106 wl_96 vdd gnd cell_6t
Xbit_r97_c106 bl_106 br_106 wl_97 vdd gnd cell_6t
Xbit_r98_c106 bl_106 br_106 wl_98 vdd gnd cell_6t
Xbit_r99_c106 bl_106 br_106 wl_99 vdd gnd cell_6t
Xbit_r100_c106 bl_106 br_106 wl_100 vdd gnd cell_6t
Xbit_r101_c106 bl_106 br_106 wl_101 vdd gnd cell_6t
Xbit_r102_c106 bl_106 br_106 wl_102 vdd gnd cell_6t
Xbit_r103_c106 bl_106 br_106 wl_103 vdd gnd cell_6t
Xbit_r104_c106 bl_106 br_106 wl_104 vdd gnd cell_6t
Xbit_r105_c106 bl_106 br_106 wl_105 vdd gnd cell_6t
Xbit_r106_c106 bl_106 br_106 wl_106 vdd gnd cell_6t
Xbit_r107_c106 bl_106 br_106 wl_107 vdd gnd cell_6t
Xbit_r108_c106 bl_106 br_106 wl_108 vdd gnd cell_6t
Xbit_r109_c106 bl_106 br_106 wl_109 vdd gnd cell_6t
Xbit_r110_c106 bl_106 br_106 wl_110 vdd gnd cell_6t
Xbit_r111_c106 bl_106 br_106 wl_111 vdd gnd cell_6t
Xbit_r112_c106 bl_106 br_106 wl_112 vdd gnd cell_6t
Xbit_r113_c106 bl_106 br_106 wl_113 vdd gnd cell_6t
Xbit_r114_c106 bl_106 br_106 wl_114 vdd gnd cell_6t
Xbit_r115_c106 bl_106 br_106 wl_115 vdd gnd cell_6t
Xbit_r116_c106 bl_106 br_106 wl_116 vdd gnd cell_6t
Xbit_r117_c106 bl_106 br_106 wl_117 vdd gnd cell_6t
Xbit_r118_c106 bl_106 br_106 wl_118 vdd gnd cell_6t
Xbit_r119_c106 bl_106 br_106 wl_119 vdd gnd cell_6t
Xbit_r120_c106 bl_106 br_106 wl_120 vdd gnd cell_6t
Xbit_r121_c106 bl_106 br_106 wl_121 vdd gnd cell_6t
Xbit_r122_c106 bl_106 br_106 wl_122 vdd gnd cell_6t
Xbit_r123_c106 bl_106 br_106 wl_123 vdd gnd cell_6t
Xbit_r124_c106 bl_106 br_106 wl_124 vdd gnd cell_6t
Xbit_r125_c106 bl_106 br_106 wl_125 vdd gnd cell_6t
Xbit_r126_c106 bl_106 br_106 wl_126 vdd gnd cell_6t
Xbit_r127_c106 bl_106 br_106 wl_127 vdd gnd cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd cell_6t
Xbit_r1_c107 bl_107 br_107 wl_1 vdd gnd cell_6t
Xbit_r2_c107 bl_107 br_107 wl_2 vdd gnd cell_6t
Xbit_r3_c107 bl_107 br_107 wl_3 vdd gnd cell_6t
Xbit_r4_c107 bl_107 br_107 wl_4 vdd gnd cell_6t
Xbit_r5_c107 bl_107 br_107 wl_5 vdd gnd cell_6t
Xbit_r6_c107 bl_107 br_107 wl_6 vdd gnd cell_6t
Xbit_r7_c107 bl_107 br_107 wl_7 vdd gnd cell_6t
Xbit_r8_c107 bl_107 br_107 wl_8 vdd gnd cell_6t
Xbit_r9_c107 bl_107 br_107 wl_9 vdd gnd cell_6t
Xbit_r10_c107 bl_107 br_107 wl_10 vdd gnd cell_6t
Xbit_r11_c107 bl_107 br_107 wl_11 vdd gnd cell_6t
Xbit_r12_c107 bl_107 br_107 wl_12 vdd gnd cell_6t
Xbit_r13_c107 bl_107 br_107 wl_13 vdd gnd cell_6t
Xbit_r14_c107 bl_107 br_107 wl_14 vdd gnd cell_6t
Xbit_r15_c107 bl_107 br_107 wl_15 vdd gnd cell_6t
Xbit_r16_c107 bl_107 br_107 wl_16 vdd gnd cell_6t
Xbit_r17_c107 bl_107 br_107 wl_17 vdd gnd cell_6t
Xbit_r18_c107 bl_107 br_107 wl_18 vdd gnd cell_6t
Xbit_r19_c107 bl_107 br_107 wl_19 vdd gnd cell_6t
Xbit_r20_c107 bl_107 br_107 wl_20 vdd gnd cell_6t
Xbit_r21_c107 bl_107 br_107 wl_21 vdd gnd cell_6t
Xbit_r22_c107 bl_107 br_107 wl_22 vdd gnd cell_6t
Xbit_r23_c107 bl_107 br_107 wl_23 vdd gnd cell_6t
Xbit_r24_c107 bl_107 br_107 wl_24 vdd gnd cell_6t
Xbit_r25_c107 bl_107 br_107 wl_25 vdd gnd cell_6t
Xbit_r26_c107 bl_107 br_107 wl_26 vdd gnd cell_6t
Xbit_r27_c107 bl_107 br_107 wl_27 vdd gnd cell_6t
Xbit_r28_c107 bl_107 br_107 wl_28 vdd gnd cell_6t
Xbit_r29_c107 bl_107 br_107 wl_29 vdd gnd cell_6t
Xbit_r30_c107 bl_107 br_107 wl_30 vdd gnd cell_6t
Xbit_r31_c107 bl_107 br_107 wl_31 vdd gnd cell_6t
Xbit_r32_c107 bl_107 br_107 wl_32 vdd gnd cell_6t
Xbit_r33_c107 bl_107 br_107 wl_33 vdd gnd cell_6t
Xbit_r34_c107 bl_107 br_107 wl_34 vdd gnd cell_6t
Xbit_r35_c107 bl_107 br_107 wl_35 vdd gnd cell_6t
Xbit_r36_c107 bl_107 br_107 wl_36 vdd gnd cell_6t
Xbit_r37_c107 bl_107 br_107 wl_37 vdd gnd cell_6t
Xbit_r38_c107 bl_107 br_107 wl_38 vdd gnd cell_6t
Xbit_r39_c107 bl_107 br_107 wl_39 vdd gnd cell_6t
Xbit_r40_c107 bl_107 br_107 wl_40 vdd gnd cell_6t
Xbit_r41_c107 bl_107 br_107 wl_41 vdd gnd cell_6t
Xbit_r42_c107 bl_107 br_107 wl_42 vdd gnd cell_6t
Xbit_r43_c107 bl_107 br_107 wl_43 vdd gnd cell_6t
Xbit_r44_c107 bl_107 br_107 wl_44 vdd gnd cell_6t
Xbit_r45_c107 bl_107 br_107 wl_45 vdd gnd cell_6t
Xbit_r46_c107 bl_107 br_107 wl_46 vdd gnd cell_6t
Xbit_r47_c107 bl_107 br_107 wl_47 vdd gnd cell_6t
Xbit_r48_c107 bl_107 br_107 wl_48 vdd gnd cell_6t
Xbit_r49_c107 bl_107 br_107 wl_49 vdd gnd cell_6t
Xbit_r50_c107 bl_107 br_107 wl_50 vdd gnd cell_6t
Xbit_r51_c107 bl_107 br_107 wl_51 vdd gnd cell_6t
Xbit_r52_c107 bl_107 br_107 wl_52 vdd gnd cell_6t
Xbit_r53_c107 bl_107 br_107 wl_53 vdd gnd cell_6t
Xbit_r54_c107 bl_107 br_107 wl_54 vdd gnd cell_6t
Xbit_r55_c107 bl_107 br_107 wl_55 vdd gnd cell_6t
Xbit_r56_c107 bl_107 br_107 wl_56 vdd gnd cell_6t
Xbit_r57_c107 bl_107 br_107 wl_57 vdd gnd cell_6t
Xbit_r58_c107 bl_107 br_107 wl_58 vdd gnd cell_6t
Xbit_r59_c107 bl_107 br_107 wl_59 vdd gnd cell_6t
Xbit_r60_c107 bl_107 br_107 wl_60 vdd gnd cell_6t
Xbit_r61_c107 bl_107 br_107 wl_61 vdd gnd cell_6t
Xbit_r62_c107 bl_107 br_107 wl_62 vdd gnd cell_6t
Xbit_r63_c107 bl_107 br_107 wl_63 vdd gnd cell_6t
Xbit_r64_c107 bl_107 br_107 wl_64 vdd gnd cell_6t
Xbit_r65_c107 bl_107 br_107 wl_65 vdd gnd cell_6t
Xbit_r66_c107 bl_107 br_107 wl_66 vdd gnd cell_6t
Xbit_r67_c107 bl_107 br_107 wl_67 vdd gnd cell_6t
Xbit_r68_c107 bl_107 br_107 wl_68 vdd gnd cell_6t
Xbit_r69_c107 bl_107 br_107 wl_69 vdd gnd cell_6t
Xbit_r70_c107 bl_107 br_107 wl_70 vdd gnd cell_6t
Xbit_r71_c107 bl_107 br_107 wl_71 vdd gnd cell_6t
Xbit_r72_c107 bl_107 br_107 wl_72 vdd gnd cell_6t
Xbit_r73_c107 bl_107 br_107 wl_73 vdd gnd cell_6t
Xbit_r74_c107 bl_107 br_107 wl_74 vdd gnd cell_6t
Xbit_r75_c107 bl_107 br_107 wl_75 vdd gnd cell_6t
Xbit_r76_c107 bl_107 br_107 wl_76 vdd gnd cell_6t
Xbit_r77_c107 bl_107 br_107 wl_77 vdd gnd cell_6t
Xbit_r78_c107 bl_107 br_107 wl_78 vdd gnd cell_6t
Xbit_r79_c107 bl_107 br_107 wl_79 vdd gnd cell_6t
Xbit_r80_c107 bl_107 br_107 wl_80 vdd gnd cell_6t
Xbit_r81_c107 bl_107 br_107 wl_81 vdd gnd cell_6t
Xbit_r82_c107 bl_107 br_107 wl_82 vdd gnd cell_6t
Xbit_r83_c107 bl_107 br_107 wl_83 vdd gnd cell_6t
Xbit_r84_c107 bl_107 br_107 wl_84 vdd gnd cell_6t
Xbit_r85_c107 bl_107 br_107 wl_85 vdd gnd cell_6t
Xbit_r86_c107 bl_107 br_107 wl_86 vdd gnd cell_6t
Xbit_r87_c107 bl_107 br_107 wl_87 vdd gnd cell_6t
Xbit_r88_c107 bl_107 br_107 wl_88 vdd gnd cell_6t
Xbit_r89_c107 bl_107 br_107 wl_89 vdd gnd cell_6t
Xbit_r90_c107 bl_107 br_107 wl_90 vdd gnd cell_6t
Xbit_r91_c107 bl_107 br_107 wl_91 vdd gnd cell_6t
Xbit_r92_c107 bl_107 br_107 wl_92 vdd gnd cell_6t
Xbit_r93_c107 bl_107 br_107 wl_93 vdd gnd cell_6t
Xbit_r94_c107 bl_107 br_107 wl_94 vdd gnd cell_6t
Xbit_r95_c107 bl_107 br_107 wl_95 vdd gnd cell_6t
Xbit_r96_c107 bl_107 br_107 wl_96 vdd gnd cell_6t
Xbit_r97_c107 bl_107 br_107 wl_97 vdd gnd cell_6t
Xbit_r98_c107 bl_107 br_107 wl_98 vdd gnd cell_6t
Xbit_r99_c107 bl_107 br_107 wl_99 vdd gnd cell_6t
Xbit_r100_c107 bl_107 br_107 wl_100 vdd gnd cell_6t
Xbit_r101_c107 bl_107 br_107 wl_101 vdd gnd cell_6t
Xbit_r102_c107 bl_107 br_107 wl_102 vdd gnd cell_6t
Xbit_r103_c107 bl_107 br_107 wl_103 vdd gnd cell_6t
Xbit_r104_c107 bl_107 br_107 wl_104 vdd gnd cell_6t
Xbit_r105_c107 bl_107 br_107 wl_105 vdd gnd cell_6t
Xbit_r106_c107 bl_107 br_107 wl_106 vdd gnd cell_6t
Xbit_r107_c107 bl_107 br_107 wl_107 vdd gnd cell_6t
Xbit_r108_c107 bl_107 br_107 wl_108 vdd gnd cell_6t
Xbit_r109_c107 bl_107 br_107 wl_109 vdd gnd cell_6t
Xbit_r110_c107 bl_107 br_107 wl_110 vdd gnd cell_6t
Xbit_r111_c107 bl_107 br_107 wl_111 vdd gnd cell_6t
Xbit_r112_c107 bl_107 br_107 wl_112 vdd gnd cell_6t
Xbit_r113_c107 bl_107 br_107 wl_113 vdd gnd cell_6t
Xbit_r114_c107 bl_107 br_107 wl_114 vdd gnd cell_6t
Xbit_r115_c107 bl_107 br_107 wl_115 vdd gnd cell_6t
Xbit_r116_c107 bl_107 br_107 wl_116 vdd gnd cell_6t
Xbit_r117_c107 bl_107 br_107 wl_117 vdd gnd cell_6t
Xbit_r118_c107 bl_107 br_107 wl_118 vdd gnd cell_6t
Xbit_r119_c107 bl_107 br_107 wl_119 vdd gnd cell_6t
Xbit_r120_c107 bl_107 br_107 wl_120 vdd gnd cell_6t
Xbit_r121_c107 bl_107 br_107 wl_121 vdd gnd cell_6t
Xbit_r122_c107 bl_107 br_107 wl_122 vdd gnd cell_6t
Xbit_r123_c107 bl_107 br_107 wl_123 vdd gnd cell_6t
Xbit_r124_c107 bl_107 br_107 wl_124 vdd gnd cell_6t
Xbit_r125_c107 bl_107 br_107 wl_125 vdd gnd cell_6t
Xbit_r126_c107 bl_107 br_107 wl_126 vdd gnd cell_6t
Xbit_r127_c107 bl_107 br_107 wl_127 vdd gnd cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd cell_6t
Xbit_r1_c108 bl_108 br_108 wl_1 vdd gnd cell_6t
Xbit_r2_c108 bl_108 br_108 wl_2 vdd gnd cell_6t
Xbit_r3_c108 bl_108 br_108 wl_3 vdd gnd cell_6t
Xbit_r4_c108 bl_108 br_108 wl_4 vdd gnd cell_6t
Xbit_r5_c108 bl_108 br_108 wl_5 vdd gnd cell_6t
Xbit_r6_c108 bl_108 br_108 wl_6 vdd gnd cell_6t
Xbit_r7_c108 bl_108 br_108 wl_7 vdd gnd cell_6t
Xbit_r8_c108 bl_108 br_108 wl_8 vdd gnd cell_6t
Xbit_r9_c108 bl_108 br_108 wl_9 vdd gnd cell_6t
Xbit_r10_c108 bl_108 br_108 wl_10 vdd gnd cell_6t
Xbit_r11_c108 bl_108 br_108 wl_11 vdd gnd cell_6t
Xbit_r12_c108 bl_108 br_108 wl_12 vdd gnd cell_6t
Xbit_r13_c108 bl_108 br_108 wl_13 vdd gnd cell_6t
Xbit_r14_c108 bl_108 br_108 wl_14 vdd gnd cell_6t
Xbit_r15_c108 bl_108 br_108 wl_15 vdd gnd cell_6t
Xbit_r16_c108 bl_108 br_108 wl_16 vdd gnd cell_6t
Xbit_r17_c108 bl_108 br_108 wl_17 vdd gnd cell_6t
Xbit_r18_c108 bl_108 br_108 wl_18 vdd gnd cell_6t
Xbit_r19_c108 bl_108 br_108 wl_19 vdd gnd cell_6t
Xbit_r20_c108 bl_108 br_108 wl_20 vdd gnd cell_6t
Xbit_r21_c108 bl_108 br_108 wl_21 vdd gnd cell_6t
Xbit_r22_c108 bl_108 br_108 wl_22 vdd gnd cell_6t
Xbit_r23_c108 bl_108 br_108 wl_23 vdd gnd cell_6t
Xbit_r24_c108 bl_108 br_108 wl_24 vdd gnd cell_6t
Xbit_r25_c108 bl_108 br_108 wl_25 vdd gnd cell_6t
Xbit_r26_c108 bl_108 br_108 wl_26 vdd gnd cell_6t
Xbit_r27_c108 bl_108 br_108 wl_27 vdd gnd cell_6t
Xbit_r28_c108 bl_108 br_108 wl_28 vdd gnd cell_6t
Xbit_r29_c108 bl_108 br_108 wl_29 vdd gnd cell_6t
Xbit_r30_c108 bl_108 br_108 wl_30 vdd gnd cell_6t
Xbit_r31_c108 bl_108 br_108 wl_31 vdd gnd cell_6t
Xbit_r32_c108 bl_108 br_108 wl_32 vdd gnd cell_6t
Xbit_r33_c108 bl_108 br_108 wl_33 vdd gnd cell_6t
Xbit_r34_c108 bl_108 br_108 wl_34 vdd gnd cell_6t
Xbit_r35_c108 bl_108 br_108 wl_35 vdd gnd cell_6t
Xbit_r36_c108 bl_108 br_108 wl_36 vdd gnd cell_6t
Xbit_r37_c108 bl_108 br_108 wl_37 vdd gnd cell_6t
Xbit_r38_c108 bl_108 br_108 wl_38 vdd gnd cell_6t
Xbit_r39_c108 bl_108 br_108 wl_39 vdd gnd cell_6t
Xbit_r40_c108 bl_108 br_108 wl_40 vdd gnd cell_6t
Xbit_r41_c108 bl_108 br_108 wl_41 vdd gnd cell_6t
Xbit_r42_c108 bl_108 br_108 wl_42 vdd gnd cell_6t
Xbit_r43_c108 bl_108 br_108 wl_43 vdd gnd cell_6t
Xbit_r44_c108 bl_108 br_108 wl_44 vdd gnd cell_6t
Xbit_r45_c108 bl_108 br_108 wl_45 vdd gnd cell_6t
Xbit_r46_c108 bl_108 br_108 wl_46 vdd gnd cell_6t
Xbit_r47_c108 bl_108 br_108 wl_47 vdd gnd cell_6t
Xbit_r48_c108 bl_108 br_108 wl_48 vdd gnd cell_6t
Xbit_r49_c108 bl_108 br_108 wl_49 vdd gnd cell_6t
Xbit_r50_c108 bl_108 br_108 wl_50 vdd gnd cell_6t
Xbit_r51_c108 bl_108 br_108 wl_51 vdd gnd cell_6t
Xbit_r52_c108 bl_108 br_108 wl_52 vdd gnd cell_6t
Xbit_r53_c108 bl_108 br_108 wl_53 vdd gnd cell_6t
Xbit_r54_c108 bl_108 br_108 wl_54 vdd gnd cell_6t
Xbit_r55_c108 bl_108 br_108 wl_55 vdd gnd cell_6t
Xbit_r56_c108 bl_108 br_108 wl_56 vdd gnd cell_6t
Xbit_r57_c108 bl_108 br_108 wl_57 vdd gnd cell_6t
Xbit_r58_c108 bl_108 br_108 wl_58 vdd gnd cell_6t
Xbit_r59_c108 bl_108 br_108 wl_59 vdd gnd cell_6t
Xbit_r60_c108 bl_108 br_108 wl_60 vdd gnd cell_6t
Xbit_r61_c108 bl_108 br_108 wl_61 vdd gnd cell_6t
Xbit_r62_c108 bl_108 br_108 wl_62 vdd gnd cell_6t
Xbit_r63_c108 bl_108 br_108 wl_63 vdd gnd cell_6t
Xbit_r64_c108 bl_108 br_108 wl_64 vdd gnd cell_6t
Xbit_r65_c108 bl_108 br_108 wl_65 vdd gnd cell_6t
Xbit_r66_c108 bl_108 br_108 wl_66 vdd gnd cell_6t
Xbit_r67_c108 bl_108 br_108 wl_67 vdd gnd cell_6t
Xbit_r68_c108 bl_108 br_108 wl_68 vdd gnd cell_6t
Xbit_r69_c108 bl_108 br_108 wl_69 vdd gnd cell_6t
Xbit_r70_c108 bl_108 br_108 wl_70 vdd gnd cell_6t
Xbit_r71_c108 bl_108 br_108 wl_71 vdd gnd cell_6t
Xbit_r72_c108 bl_108 br_108 wl_72 vdd gnd cell_6t
Xbit_r73_c108 bl_108 br_108 wl_73 vdd gnd cell_6t
Xbit_r74_c108 bl_108 br_108 wl_74 vdd gnd cell_6t
Xbit_r75_c108 bl_108 br_108 wl_75 vdd gnd cell_6t
Xbit_r76_c108 bl_108 br_108 wl_76 vdd gnd cell_6t
Xbit_r77_c108 bl_108 br_108 wl_77 vdd gnd cell_6t
Xbit_r78_c108 bl_108 br_108 wl_78 vdd gnd cell_6t
Xbit_r79_c108 bl_108 br_108 wl_79 vdd gnd cell_6t
Xbit_r80_c108 bl_108 br_108 wl_80 vdd gnd cell_6t
Xbit_r81_c108 bl_108 br_108 wl_81 vdd gnd cell_6t
Xbit_r82_c108 bl_108 br_108 wl_82 vdd gnd cell_6t
Xbit_r83_c108 bl_108 br_108 wl_83 vdd gnd cell_6t
Xbit_r84_c108 bl_108 br_108 wl_84 vdd gnd cell_6t
Xbit_r85_c108 bl_108 br_108 wl_85 vdd gnd cell_6t
Xbit_r86_c108 bl_108 br_108 wl_86 vdd gnd cell_6t
Xbit_r87_c108 bl_108 br_108 wl_87 vdd gnd cell_6t
Xbit_r88_c108 bl_108 br_108 wl_88 vdd gnd cell_6t
Xbit_r89_c108 bl_108 br_108 wl_89 vdd gnd cell_6t
Xbit_r90_c108 bl_108 br_108 wl_90 vdd gnd cell_6t
Xbit_r91_c108 bl_108 br_108 wl_91 vdd gnd cell_6t
Xbit_r92_c108 bl_108 br_108 wl_92 vdd gnd cell_6t
Xbit_r93_c108 bl_108 br_108 wl_93 vdd gnd cell_6t
Xbit_r94_c108 bl_108 br_108 wl_94 vdd gnd cell_6t
Xbit_r95_c108 bl_108 br_108 wl_95 vdd gnd cell_6t
Xbit_r96_c108 bl_108 br_108 wl_96 vdd gnd cell_6t
Xbit_r97_c108 bl_108 br_108 wl_97 vdd gnd cell_6t
Xbit_r98_c108 bl_108 br_108 wl_98 vdd gnd cell_6t
Xbit_r99_c108 bl_108 br_108 wl_99 vdd gnd cell_6t
Xbit_r100_c108 bl_108 br_108 wl_100 vdd gnd cell_6t
Xbit_r101_c108 bl_108 br_108 wl_101 vdd gnd cell_6t
Xbit_r102_c108 bl_108 br_108 wl_102 vdd gnd cell_6t
Xbit_r103_c108 bl_108 br_108 wl_103 vdd gnd cell_6t
Xbit_r104_c108 bl_108 br_108 wl_104 vdd gnd cell_6t
Xbit_r105_c108 bl_108 br_108 wl_105 vdd gnd cell_6t
Xbit_r106_c108 bl_108 br_108 wl_106 vdd gnd cell_6t
Xbit_r107_c108 bl_108 br_108 wl_107 vdd gnd cell_6t
Xbit_r108_c108 bl_108 br_108 wl_108 vdd gnd cell_6t
Xbit_r109_c108 bl_108 br_108 wl_109 vdd gnd cell_6t
Xbit_r110_c108 bl_108 br_108 wl_110 vdd gnd cell_6t
Xbit_r111_c108 bl_108 br_108 wl_111 vdd gnd cell_6t
Xbit_r112_c108 bl_108 br_108 wl_112 vdd gnd cell_6t
Xbit_r113_c108 bl_108 br_108 wl_113 vdd gnd cell_6t
Xbit_r114_c108 bl_108 br_108 wl_114 vdd gnd cell_6t
Xbit_r115_c108 bl_108 br_108 wl_115 vdd gnd cell_6t
Xbit_r116_c108 bl_108 br_108 wl_116 vdd gnd cell_6t
Xbit_r117_c108 bl_108 br_108 wl_117 vdd gnd cell_6t
Xbit_r118_c108 bl_108 br_108 wl_118 vdd gnd cell_6t
Xbit_r119_c108 bl_108 br_108 wl_119 vdd gnd cell_6t
Xbit_r120_c108 bl_108 br_108 wl_120 vdd gnd cell_6t
Xbit_r121_c108 bl_108 br_108 wl_121 vdd gnd cell_6t
Xbit_r122_c108 bl_108 br_108 wl_122 vdd gnd cell_6t
Xbit_r123_c108 bl_108 br_108 wl_123 vdd gnd cell_6t
Xbit_r124_c108 bl_108 br_108 wl_124 vdd gnd cell_6t
Xbit_r125_c108 bl_108 br_108 wl_125 vdd gnd cell_6t
Xbit_r126_c108 bl_108 br_108 wl_126 vdd gnd cell_6t
Xbit_r127_c108 bl_108 br_108 wl_127 vdd gnd cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd cell_6t
Xbit_r1_c109 bl_109 br_109 wl_1 vdd gnd cell_6t
Xbit_r2_c109 bl_109 br_109 wl_2 vdd gnd cell_6t
Xbit_r3_c109 bl_109 br_109 wl_3 vdd gnd cell_6t
Xbit_r4_c109 bl_109 br_109 wl_4 vdd gnd cell_6t
Xbit_r5_c109 bl_109 br_109 wl_5 vdd gnd cell_6t
Xbit_r6_c109 bl_109 br_109 wl_6 vdd gnd cell_6t
Xbit_r7_c109 bl_109 br_109 wl_7 vdd gnd cell_6t
Xbit_r8_c109 bl_109 br_109 wl_8 vdd gnd cell_6t
Xbit_r9_c109 bl_109 br_109 wl_9 vdd gnd cell_6t
Xbit_r10_c109 bl_109 br_109 wl_10 vdd gnd cell_6t
Xbit_r11_c109 bl_109 br_109 wl_11 vdd gnd cell_6t
Xbit_r12_c109 bl_109 br_109 wl_12 vdd gnd cell_6t
Xbit_r13_c109 bl_109 br_109 wl_13 vdd gnd cell_6t
Xbit_r14_c109 bl_109 br_109 wl_14 vdd gnd cell_6t
Xbit_r15_c109 bl_109 br_109 wl_15 vdd gnd cell_6t
Xbit_r16_c109 bl_109 br_109 wl_16 vdd gnd cell_6t
Xbit_r17_c109 bl_109 br_109 wl_17 vdd gnd cell_6t
Xbit_r18_c109 bl_109 br_109 wl_18 vdd gnd cell_6t
Xbit_r19_c109 bl_109 br_109 wl_19 vdd gnd cell_6t
Xbit_r20_c109 bl_109 br_109 wl_20 vdd gnd cell_6t
Xbit_r21_c109 bl_109 br_109 wl_21 vdd gnd cell_6t
Xbit_r22_c109 bl_109 br_109 wl_22 vdd gnd cell_6t
Xbit_r23_c109 bl_109 br_109 wl_23 vdd gnd cell_6t
Xbit_r24_c109 bl_109 br_109 wl_24 vdd gnd cell_6t
Xbit_r25_c109 bl_109 br_109 wl_25 vdd gnd cell_6t
Xbit_r26_c109 bl_109 br_109 wl_26 vdd gnd cell_6t
Xbit_r27_c109 bl_109 br_109 wl_27 vdd gnd cell_6t
Xbit_r28_c109 bl_109 br_109 wl_28 vdd gnd cell_6t
Xbit_r29_c109 bl_109 br_109 wl_29 vdd gnd cell_6t
Xbit_r30_c109 bl_109 br_109 wl_30 vdd gnd cell_6t
Xbit_r31_c109 bl_109 br_109 wl_31 vdd gnd cell_6t
Xbit_r32_c109 bl_109 br_109 wl_32 vdd gnd cell_6t
Xbit_r33_c109 bl_109 br_109 wl_33 vdd gnd cell_6t
Xbit_r34_c109 bl_109 br_109 wl_34 vdd gnd cell_6t
Xbit_r35_c109 bl_109 br_109 wl_35 vdd gnd cell_6t
Xbit_r36_c109 bl_109 br_109 wl_36 vdd gnd cell_6t
Xbit_r37_c109 bl_109 br_109 wl_37 vdd gnd cell_6t
Xbit_r38_c109 bl_109 br_109 wl_38 vdd gnd cell_6t
Xbit_r39_c109 bl_109 br_109 wl_39 vdd gnd cell_6t
Xbit_r40_c109 bl_109 br_109 wl_40 vdd gnd cell_6t
Xbit_r41_c109 bl_109 br_109 wl_41 vdd gnd cell_6t
Xbit_r42_c109 bl_109 br_109 wl_42 vdd gnd cell_6t
Xbit_r43_c109 bl_109 br_109 wl_43 vdd gnd cell_6t
Xbit_r44_c109 bl_109 br_109 wl_44 vdd gnd cell_6t
Xbit_r45_c109 bl_109 br_109 wl_45 vdd gnd cell_6t
Xbit_r46_c109 bl_109 br_109 wl_46 vdd gnd cell_6t
Xbit_r47_c109 bl_109 br_109 wl_47 vdd gnd cell_6t
Xbit_r48_c109 bl_109 br_109 wl_48 vdd gnd cell_6t
Xbit_r49_c109 bl_109 br_109 wl_49 vdd gnd cell_6t
Xbit_r50_c109 bl_109 br_109 wl_50 vdd gnd cell_6t
Xbit_r51_c109 bl_109 br_109 wl_51 vdd gnd cell_6t
Xbit_r52_c109 bl_109 br_109 wl_52 vdd gnd cell_6t
Xbit_r53_c109 bl_109 br_109 wl_53 vdd gnd cell_6t
Xbit_r54_c109 bl_109 br_109 wl_54 vdd gnd cell_6t
Xbit_r55_c109 bl_109 br_109 wl_55 vdd gnd cell_6t
Xbit_r56_c109 bl_109 br_109 wl_56 vdd gnd cell_6t
Xbit_r57_c109 bl_109 br_109 wl_57 vdd gnd cell_6t
Xbit_r58_c109 bl_109 br_109 wl_58 vdd gnd cell_6t
Xbit_r59_c109 bl_109 br_109 wl_59 vdd gnd cell_6t
Xbit_r60_c109 bl_109 br_109 wl_60 vdd gnd cell_6t
Xbit_r61_c109 bl_109 br_109 wl_61 vdd gnd cell_6t
Xbit_r62_c109 bl_109 br_109 wl_62 vdd gnd cell_6t
Xbit_r63_c109 bl_109 br_109 wl_63 vdd gnd cell_6t
Xbit_r64_c109 bl_109 br_109 wl_64 vdd gnd cell_6t
Xbit_r65_c109 bl_109 br_109 wl_65 vdd gnd cell_6t
Xbit_r66_c109 bl_109 br_109 wl_66 vdd gnd cell_6t
Xbit_r67_c109 bl_109 br_109 wl_67 vdd gnd cell_6t
Xbit_r68_c109 bl_109 br_109 wl_68 vdd gnd cell_6t
Xbit_r69_c109 bl_109 br_109 wl_69 vdd gnd cell_6t
Xbit_r70_c109 bl_109 br_109 wl_70 vdd gnd cell_6t
Xbit_r71_c109 bl_109 br_109 wl_71 vdd gnd cell_6t
Xbit_r72_c109 bl_109 br_109 wl_72 vdd gnd cell_6t
Xbit_r73_c109 bl_109 br_109 wl_73 vdd gnd cell_6t
Xbit_r74_c109 bl_109 br_109 wl_74 vdd gnd cell_6t
Xbit_r75_c109 bl_109 br_109 wl_75 vdd gnd cell_6t
Xbit_r76_c109 bl_109 br_109 wl_76 vdd gnd cell_6t
Xbit_r77_c109 bl_109 br_109 wl_77 vdd gnd cell_6t
Xbit_r78_c109 bl_109 br_109 wl_78 vdd gnd cell_6t
Xbit_r79_c109 bl_109 br_109 wl_79 vdd gnd cell_6t
Xbit_r80_c109 bl_109 br_109 wl_80 vdd gnd cell_6t
Xbit_r81_c109 bl_109 br_109 wl_81 vdd gnd cell_6t
Xbit_r82_c109 bl_109 br_109 wl_82 vdd gnd cell_6t
Xbit_r83_c109 bl_109 br_109 wl_83 vdd gnd cell_6t
Xbit_r84_c109 bl_109 br_109 wl_84 vdd gnd cell_6t
Xbit_r85_c109 bl_109 br_109 wl_85 vdd gnd cell_6t
Xbit_r86_c109 bl_109 br_109 wl_86 vdd gnd cell_6t
Xbit_r87_c109 bl_109 br_109 wl_87 vdd gnd cell_6t
Xbit_r88_c109 bl_109 br_109 wl_88 vdd gnd cell_6t
Xbit_r89_c109 bl_109 br_109 wl_89 vdd gnd cell_6t
Xbit_r90_c109 bl_109 br_109 wl_90 vdd gnd cell_6t
Xbit_r91_c109 bl_109 br_109 wl_91 vdd gnd cell_6t
Xbit_r92_c109 bl_109 br_109 wl_92 vdd gnd cell_6t
Xbit_r93_c109 bl_109 br_109 wl_93 vdd gnd cell_6t
Xbit_r94_c109 bl_109 br_109 wl_94 vdd gnd cell_6t
Xbit_r95_c109 bl_109 br_109 wl_95 vdd gnd cell_6t
Xbit_r96_c109 bl_109 br_109 wl_96 vdd gnd cell_6t
Xbit_r97_c109 bl_109 br_109 wl_97 vdd gnd cell_6t
Xbit_r98_c109 bl_109 br_109 wl_98 vdd gnd cell_6t
Xbit_r99_c109 bl_109 br_109 wl_99 vdd gnd cell_6t
Xbit_r100_c109 bl_109 br_109 wl_100 vdd gnd cell_6t
Xbit_r101_c109 bl_109 br_109 wl_101 vdd gnd cell_6t
Xbit_r102_c109 bl_109 br_109 wl_102 vdd gnd cell_6t
Xbit_r103_c109 bl_109 br_109 wl_103 vdd gnd cell_6t
Xbit_r104_c109 bl_109 br_109 wl_104 vdd gnd cell_6t
Xbit_r105_c109 bl_109 br_109 wl_105 vdd gnd cell_6t
Xbit_r106_c109 bl_109 br_109 wl_106 vdd gnd cell_6t
Xbit_r107_c109 bl_109 br_109 wl_107 vdd gnd cell_6t
Xbit_r108_c109 bl_109 br_109 wl_108 vdd gnd cell_6t
Xbit_r109_c109 bl_109 br_109 wl_109 vdd gnd cell_6t
Xbit_r110_c109 bl_109 br_109 wl_110 vdd gnd cell_6t
Xbit_r111_c109 bl_109 br_109 wl_111 vdd gnd cell_6t
Xbit_r112_c109 bl_109 br_109 wl_112 vdd gnd cell_6t
Xbit_r113_c109 bl_109 br_109 wl_113 vdd gnd cell_6t
Xbit_r114_c109 bl_109 br_109 wl_114 vdd gnd cell_6t
Xbit_r115_c109 bl_109 br_109 wl_115 vdd gnd cell_6t
Xbit_r116_c109 bl_109 br_109 wl_116 vdd gnd cell_6t
Xbit_r117_c109 bl_109 br_109 wl_117 vdd gnd cell_6t
Xbit_r118_c109 bl_109 br_109 wl_118 vdd gnd cell_6t
Xbit_r119_c109 bl_109 br_109 wl_119 vdd gnd cell_6t
Xbit_r120_c109 bl_109 br_109 wl_120 vdd gnd cell_6t
Xbit_r121_c109 bl_109 br_109 wl_121 vdd gnd cell_6t
Xbit_r122_c109 bl_109 br_109 wl_122 vdd gnd cell_6t
Xbit_r123_c109 bl_109 br_109 wl_123 vdd gnd cell_6t
Xbit_r124_c109 bl_109 br_109 wl_124 vdd gnd cell_6t
Xbit_r125_c109 bl_109 br_109 wl_125 vdd gnd cell_6t
Xbit_r126_c109 bl_109 br_109 wl_126 vdd gnd cell_6t
Xbit_r127_c109 bl_109 br_109 wl_127 vdd gnd cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd cell_6t
Xbit_r1_c110 bl_110 br_110 wl_1 vdd gnd cell_6t
Xbit_r2_c110 bl_110 br_110 wl_2 vdd gnd cell_6t
Xbit_r3_c110 bl_110 br_110 wl_3 vdd gnd cell_6t
Xbit_r4_c110 bl_110 br_110 wl_4 vdd gnd cell_6t
Xbit_r5_c110 bl_110 br_110 wl_5 vdd gnd cell_6t
Xbit_r6_c110 bl_110 br_110 wl_6 vdd gnd cell_6t
Xbit_r7_c110 bl_110 br_110 wl_7 vdd gnd cell_6t
Xbit_r8_c110 bl_110 br_110 wl_8 vdd gnd cell_6t
Xbit_r9_c110 bl_110 br_110 wl_9 vdd gnd cell_6t
Xbit_r10_c110 bl_110 br_110 wl_10 vdd gnd cell_6t
Xbit_r11_c110 bl_110 br_110 wl_11 vdd gnd cell_6t
Xbit_r12_c110 bl_110 br_110 wl_12 vdd gnd cell_6t
Xbit_r13_c110 bl_110 br_110 wl_13 vdd gnd cell_6t
Xbit_r14_c110 bl_110 br_110 wl_14 vdd gnd cell_6t
Xbit_r15_c110 bl_110 br_110 wl_15 vdd gnd cell_6t
Xbit_r16_c110 bl_110 br_110 wl_16 vdd gnd cell_6t
Xbit_r17_c110 bl_110 br_110 wl_17 vdd gnd cell_6t
Xbit_r18_c110 bl_110 br_110 wl_18 vdd gnd cell_6t
Xbit_r19_c110 bl_110 br_110 wl_19 vdd gnd cell_6t
Xbit_r20_c110 bl_110 br_110 wl_20 vdd gnd cell_6t
Xbit_r21_c110 bl_110 br_110 wl_21 vdd gnd cell_6t
Xbit_r22_c110 bl_110 br_110 wl_22 vdd gnd cell_6t
Xbit_r23_c110 bl_110 br_110 wl_23 vdd gnd cell_6t
Xbit_r24_c110 bl_110 br_110 wl_24 vdd gnd cell_6t
Xbit_r25_c110 bl_110 br_110 wl_25 vdd gnd cell_6t
Xbit_r26_c110 bl_110 br_110 wl_26 vdd gnd cell_6t
Xbit_r27_c110 bl_110 br_110 wl_27 vdd gnd cell_6t
Xbit_r28_c110 bl_110 br_110 wl_28 vdd gnd cell_6t
Xbit_r29_c110 bl_110 br_110 wl_29 vdd gnd cell_6t
Xbit_r30_c110 bl_110 br_110 wl_30 vdd gnd cell_6t
Xbit_r31_c110 bl_110 br_110 wl_31 vdd gnd cell_6t
Xbit_r32_c110 bl_110 br_110 wl_32 vdd gnd cell_6t
Xbit_r33_c110 bl_110 br_110 wl_33 vdd gnd cell_6t
Xbit_r34_c110 bl_110 br_110 wl_34 vdd gnd cell_6t
Xbit_r35_c110 bl_110 br_110 wl_35 vdd gnd cell_6t
Xbit_r36_c110 bl_110 br_110 wl_36 vdd gnd cell_6t
Xbit_r37_c110 bl_110 br_110 wl_37 vdd gnd cell_6t
Xbit_r38_c110 bl_110 br_110 wl_38 vdd gnd cell_6t
Xbit_r39_c110 bl_110 br_110 wl_39 vdd gnd cell_6t
Xbit_r40_c110 bl_110 br_110 wl_40 vdd gnd cell_6t
Xbit_r41_c110 bl_110 br_110 wl_41 vdd gnd cell_6t
Xbit_r42_c110 bl_110 br_110 wl_42 vdd gnd cell_6t
Xbit_r43_c110 bl_110 br_110 wl_43 vdd gnd cell_6t
Xbit_r44_c110 bl_110 br_110 wl_44 vdd gnd cell_6t
Xbit_r45_c110 bl_110 br_110 wl_45 vdd gnd cell_6t
Xbit_r46_c110 bl_110 br_110 wl_46 vdd gnd cell_6t
Xbit_r47_c110 bl_110 br_110 wl_47 vdd gnd cell_6t
Xbit_r48_c110 bl_110 br_110 wl_48 vdd gnd cell_6t
Xbit_r49_c110 bl_110 br_110 wl_49 vdd gnd cell_6t
Xbit_r50_c110 bl_110 br_110 wl_50 vdd gnd cell_6t
Xbit_r51_c110 bl_110 br_110 wl_51 vdd gnd cell_6t
Xbit_r52_c110 bl_110 br_110 wl_52 vdd gnd cell_6t
Xbit_r53_c110 bl_110 br_110 wl_53 vdd gnd cell_6t
Xbit_r54_c110 bl_110 br_110 wl_54 vdd gnd cell_6t
Xbit_r55_c110 bl_110 br_110 wl_55 vdd gnd cell_6t
Xbit_r56_c110 bl_110 br_110 wl_56 vdd gnd cell_6t
Xbit_r57_c110 bl_110 br_110 wl_57 vdd gnd cell_6t
Xbit_r58_c110 bl_110 br_110 wl_58 vdd gnd cell_6t
Xbit_r59_c110 bl_110 br_110 wl_59 vdd gnd cell_6t
Xbit_r60_c110 bl_110 br_110 wl_60 vdd gnd cell_6t
Xbit_r61_c110 bl_110 br_110 wl_61 vdd gnd cell_6t
Xbit_r62_c110 bl_110 br_110 wl_62 vdd gnd cell_6t
Xbit_r63_c110 bl_110 br_110 wl_63 vdd gnd cell_6t
Xbit_r64_c110 bl_110 br_110 wl_64 vdd gnd cell_6t
Xbit_r65_c110 bl_110 br_110 wl_65 vdd gnd cell_6t
Xbit_r66_c110 bl_110 br_110 wl_66 vdd gnd cell_6t
Xbit_r67_c110 bl_110 br_110 wl_67 vdd gnd cell_6t
Xbit_r68_c110 bl_110 br_110 wl_68 vdd gnd cell_6t
Xbit_r69_c110 bl_110 br_110 wl_69 vdd gnd cell_6t
Xbit_r70_c110 bl_110 br_110 wl_70 vdd gnd cell_6t
Xbit_r71_c110 bl_110 br_110 wl_71 vdd gnd cell_6t
Xbit_r72_c110 bl_110 br_110 wl_72 vdd gnd cell_6t
Xbit_r73_c110 bl_110 br_110 wl_73 vdd gnd cell_6t
Xbit_r74_c110 bl_110 br_110 wl_74 vdd gnd cell_6t
Xbit_r75_c110 bl_110 br_110 wl_75 vdd gnd cell_6t
Xbit_r76_c110 bl_110 br_110 wl_76 vdd gnd cell_6t
Xbit_r77_c110 bl_110 br_110 wl_77 vdd gnd cell_6t
Xbit_r78_c110 bl_110 br_110 wl_78 vdd gnd cell_6t
Xbit_r79_c110 bl_110 br_110 wl_79 vdd gnd cell_6t
Xbit_r80_c110 bl_110 br_110 wl_80 vdd gnd cell_6t
Xbit_r81_c110 bl_110 br_110 wl_81 vdd gnd cell_6t
Xbit_r82_c110 bl_110 br_110 wl_82 vdd gnd cell_6t
Xbit_r83_c110 bl_110 br_110 wl_83 vdd gnd cell_6t
Xbit_r84_c110 bl_110 br_110 wl_84 vdd gnd cell_6t
Xbit_r85_c110 bl_110 br_110 wl_85 vdd gnd cell_6t
Xbit_r86_c110 bl_110 br_110 wl_86 vdd gnd cell_6t
Xbit_r87_c110 bl_110 br_110 wl_87 vdd gnd cell_6t
Xbit_r88_c110 bl_110 br_110 wl_88 vdd gnd cell_6t
Xbit_r89_c110 bl_110 br_110 wl_89 vdd gnd cell_6t
Xbit_r90_c110 bl_110 br_110 wl_90 vdd gnd cell_6t
Xbit_r91_c110 bl_110 br_110 wl_91 vdd gnd cell_6t
Xbit_r92_c110 bl_110 br_110 wl_92 vdd gnd cell_6t
Xbit_r93_c110 bl_110 br_110 wl_93 vdd gnd cell_6t
Xbit_r94_c110 bl_110 br_110 wl_94 vdd gnd cell_6t
Xbit_r95_c110 bl_110 br_110 wl_95 vdd gnd cell_6t
Xbit_r96_c110 bl_110 br_110 wl_96 vdd gnd cell_6t
Xbit_r97_c110 bl_110 br_110 wl_97 vdd gnd cell_6t
Xbit_r98_c110 bl_110 br_110 wl_98 vdd gnd cell_6t
Xbit_r99_c110 bl_110 br_110 wl_99 vdd gnd cell_6t
Xbit_r100_c110 bl_110 br_110 wl_100 vdd gnd cell_6t
Xbit_r101_c110 bl_110 br_110 wl_101 vdd gnd cell_6t
Xbit_r102_c110 bl_110 br_110 wl_102 vdd gnd cell_6t
Xbit_r103_c110 bl_110 br_110 wl_103 vdd gnd cell_6t
Xbit_r104_c110 bl_110 br_110 wl_104 vdd gnd cell_6t
Xbit_r105_c110 bl_110 br_110 wl_105 vdd gnd cell_6t
Xbit_r106_c110 bl_110 br_110 wl_106 vdd gnd cell_6t
Xbit_r107_c110 bl_110 br_110 wl_107 vdd gnd cell_6t
Xbit_r108_c110 bl_110 br_110 wl_108 vdd gnd cell_6t
Xbit_r109_c110 bl_110 br_110 wl_109 vdd gnd cell_6t
Xbit_r110_c110 bl_110 br_110 wl_110 vdd gnd cell_6t
Xbit_r111_c110 bl_110 br_110 wl_111 vdd gnd cell_6t
Xbit_r112_c110 bl_110 br_110 wl_112 vdd gnd cell_6t
Xbit_r113_c110 bl_110 br_110 wl_113 vdd gnd cell_6t
Xbit_r114_c110 bl_110 br_110 wl_114 vdd gnd cell_6t
Xbit_r115_c110 bl_110 br_110 wl_115 vdd gnd cell_6t
Xbit_r116_c110 bl_110 br_110 wl_116 vdd gnd cell_6t
Xbit_r117_c110 bl_110 br_110 wl_117 vdd gnd cell_6t
Xbit_r118_c110 bl_110 br_110 wl_118 vdd gnd cell_6t
Xbit_r119_c110 bl_110 br_110 wl_119 vdd gnd cell_6t
Xbit_r120_c110 bl_110 br_110 wl_120 vdd gnd cell_6t
Xbit_r121_c110 bl_110 br_110 wl_121 vdd gnd cell_6t
Xbit_r122_c110 bl_110 br_110 wl_122 vdd gnd cell_6t
Xbit_r123_c110 bl_110 br_110 wl_123 vdd gnd cell_6t
Xbit_r124_c110 bl_110 br_110 wl_124 vdd gnd cell_6t
Xbit_r125_c110 bl_110 br_110 wl_125 vdd gnd cell_6t
Xbit_r126_c110 bl_110 br_110 wl_126 vdd gnd cell_6t
Xbit_r127_c110 bl_110 br_110 wl_127 vdd gnd cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd cell_6t
Xbit_r1_c111 bl_111 br_111 wl_1 vdd gnd cell_6t
Xbit_r2_c111 bl_111 br_111 wl_2 vdd gnd cell_6t
Xbit_r3_c111 bl_111 br_111 wl_3 vdd gnd cell_6t
Xbit_r4_c111 bl_111 br_111 wl_4 vdd gnd cell_6t
Xbit_r5_c111 bl_111 br_111 wl_5 vdd gnd cell_6t
Xbit_r6_c111 bl_111 br_111 wl_6 vdd gnd cell_6t
Xbit_r7_c111 bl_111 br_111 wl_7 vdd gnd cell_6t
Xbit_r8_c111 bl_111 br_111 wl_8 vdd gnd cell_6t
Xbit_r9_c111 bl_111 br_111 wl_9 vdd gnd cell_6t
Xbit_r10_c111 bl_111 br_111 wl_10 vdd gnd cell_6t
Xbit_r11_c111 bl_111 br_111 wl_11 vdd gnd cell_6t
Xbit_r12_c111 bl_111 br_111 wl_12 vdd gnd cell_6t
Xbit_r13_c111 bl_111 br_111 wl_13 vdd gnd cell_6t
Xbit_r14_c111 bl_111 br_111 wl_14 vdd gnd cell_6t
Xbit_r15_c111 bl_111 br_111 wl_15 vdd gnd cell_6t
Xbit_r16_c111 bl_111 br_111 wl_16 vdd gnd cell_6t
Xbit_r17_c111 bl_111 br_111 wl_17 vdd gnd cell_6t
Xbit_r18_c111 bl_111 br_111 wl_18 vdd gnd cell_6t
Xbit_r19_c111 bl_111 br_111 wl_19 vdd gnd cell_6t
Xbit_r20_c111 bl_111 br_111 wl_20 vdd gnd cell_6t
Xbit_r21_c111 bl_111 br_111 wl_21 vdd gnd cell_6t
Xbit_r22_c111 bl_111 br_111 wl_22 vdd gnd cell_6t
Xbit_r23_c111 bl_111 br_111 wl_23 vdd gnd cell_6t
Xbit_r24_c111 bl_111 br_111 wl_24 vdd gnd cell_6t
Xbit_r25_c111 bl_111 br_111 wl_25 vdd gnd cell_6t
Xbit_r26_c111 bl_111 br_111 wl_26 vdd gnd cell_6t
Xbit_r27_c111 bl_111 br_111 wl_27 vdd gnd cell_6t
Xbit_r28_c111 bl_111 br_111 wl_28 vdd gnd cell_6t
Xbit_r29_c111 bl_111 br_111 wl_29 vdd gnd cell_6t
Xbit_r30_c111 bl_111 br_111 wl_30 vdd gnd cell_6t
Xbit_r31_c111 bl_111 br_111 wl_31 vdd gnd cell_6t
Xbit_r32_c111 bl_111 br_111 wl_32 vdd gnd cell_6t
Xbit_r33_c111 bl_111 br_111 wl_33 vdd gnd cell_6t
Xbit_r34_c111 bl_111 br_111 wl_34 vdd gnd cell_6t
Xbit_r35_c111 bl_111 br_111 wl_35 vdd gnd cell_6t
Xbit_r36_c111 bl_111 br_111 wl_36 vdd gnd cell_6t
Xbit_r37_c111 bl_111 br_111 wl_37 vdd gnd cell_6t
Xbit_r38_c111 bl_111 br_111 wl_38 vdd gnd cell_6t
Xbit_r39_c111 bl_111 br_111 wl_39 vdd gnd cell_6t
Xbit_r40_c111 bl_111 br_111 wl_40 vdd gnd cell_6t
Xbit_r41_c111 bl_111 br_111 wl_41 vdd gnd cell_6t
Xbit_r42_c111 bl_111 br_111 wl_42 vdd gnd cell_6t
Xbit_r43_c111 bl_111 br_111 wl_43 vdd gnd cell_6t
Xbit_r44_c111 bl_111 br_111 wl_44 vdd gnd cell_6t
Xbit_r45_c111 bl_111 br_111 wl_45 vdd gnd cell_6t
Xbit_r46_c111 bl_111 br_111 wl_46 vdd gnd cell_6t
Xbit_r47_c111 bl_111 br_111 wl_47 vdd gnd cell_6t
Xbit_r48_c111 bl_111 br_111 wl_48 vdd gnd cell_6t
Xbit_r49_c111 bl_111 br_111 wl_49 vdd gnd cell_6t
Xbit_r50_c111 bl_111 br_111 wl_50 vdd gnd cell_6t
Xbit_r51_c111 bl_111 br_111 wl_51 vdd gnd cell_6t
Xbit_r52_c111 bl_111 br_111 wl_52 vdd gnd cell_6t
Xbit_r53_c111 bl_111 br_111 wl_53 vdd gnd cell_6t
Xbit_r54_c111 bl_111 br_111 wl_54 vdd gnd cell_6t
Xbit_r55_c111 bl_111 br_111 wl_55 vdd gnd cell_6t
Xbit_r56_c111 bl_111 br_111 wl_56 vdd gnd cell_6t
Xbit_r57_c111 bl_111 br_111 wl_57 vdd gnd cell_6t
Xbit_r58_c111 bl_111 br_111 wl_58 vdd gnd cell_6t
Xbit_r59_c111 bl_111 br_111 wl_59 vdd gnd cell_6t
Xbit_r60_c111 bl_111 br_111 wl_60 vdd gnd cell_6t
Xbit_r61_c111 bl_111 br_111 wl_61 vdd gnd cell_6t
Xbit_r62_c111 bl_111 br_111 wl_62 vdd gnd cell_6t
Xbit_r63_c111 bl_111 br_111 wl_63 vdd gnd cell_6t
Xbit_r64_c111 bl_111 br_111 wl_64 vdd gnd cell_6t
Xbit_r65_c111 bl_111 br_111 wl_65 vdd gnd cell_6t
Xbit_r66_c111 bl_111 br_111 wl_66 vdd gnd cell_6t
Xbit_r67_c111 bl_111 br_111 wl_67 vdd gnd cell_6t
Xbit_r68_c111 bl_111 br_111 wl_68 vdd gnd cell_6t
Xbit_r69_c111 bl_111 br_111 wl_69 vdd gnd cell_6t
Xbit_r70_c111 bl_111 br_111 wl_70 vdd gnd cell_6t
Xbit_r71_c111 bl_111 br_111 wl_71 vdd gnd cell_6t
Xbit_r72_c111 bl_111 br_111 wl_72 vdd gnd cell_6t
Xbit_r73_c111 bl_111 br_111 wl_73 vdd gnd cell_6t
Xbit_r74_c111 bl_111 br_111 wl_74 vdd gnd cell_6t
Xbit_r75_c111 bl_111 br_111 wl_75 vdd gnd cell_6t
Xbit_r76_c111 bl_111 br_111 wl_76 vdd gnd cell_6t
Xbit_r77_c111 bl_111 br_111 wl_77 vdd gnd cell_6t
Xbit_r78_c111 bl_111 br_111 wl_78 vdd gnd cell_6t
Xbit_r79_c111 bl_111 br_111 wl_79 vdd gnd cell_6t
Xbit_r80_c111 bl_111 br_111 wl_80 vdd gnd cell_6t
Xbit_r81_c111 bl_111 br_111 wl_81 vdd gnd cell_6t
Xbit_r82_c111 bl_111 br_111 wl_82 vdd gnd cell_6t
Xbit_r83_c111 bl_111 br_111 wl_83 vdd gnd cell_6t
Xbit_r84_c111 bl_111 br_111 wl_84 vdd gnd cell_6t
Xbit_r85_c111 bl_111 br_111 wl_85 vdd gnd cell_6t
Xbit_r86_c111 bl_111 br_111 wl_86 vdd gnd cell_6t
Xbit_r87_c111 bl_111 br_111 wl_87 vdd gnd cell_6t
Xbit_r88_c111 bl_111 br_111 wl_88 vdd gnd cell_6t
Xbit_r89_c111 bl_111 br_111 wl_89 vdd gnd cell_6t
Xbit_r90_c111 bl_111 br_111 wl_90 vdd gnd cell_6t
Xbit_r91_c111 bl_111 br_111 wl_91 vdd gnd cell_6t
Xbit_r92_c111 bl_111 br_111 wl_92 vdd gnd cell_6t
Xbit_r93_c111 bl_111 br_111 wl_93 vdd gnd cell_6t
Xbit_r94_c111 bl_111 br_111 wl_94 vdd gnd cell_6t
Xbit_r95_c111 bl_111 br_111 wl_95 vdd gnd cell_6t
Xbit_r96_c111 bl_111 br_111 wl_96 vdd gnd cell_6t
Xbit_r97_c111 bl_111 br_111 wl_97 vdd gnd cell_6t
Xbit_r98_c111 bl_111 br_111 wl_98 vdd gnd cell_6t
Xbit_r99_c111 bl_111 br_111 wl_99 vdd gnd cell_6t
Xbit_r100_c111 bl_111 br_111 wl_100 vdd gnd cell_6t
Xbit_r101_c111 bl_111 br_111 wl_101 vdd gnd cell_6t
Xbit_r102_c111 bl_111 br_111 wl_102 vdd gnd cell_6t
Xbit_r103_c111 bl_111 br_111 wl_103 vdd gnd cell_6t
Xbit_r104_c111 bl_111 br_111 wl_104 vdd gnd cell_6t
Xbit_r105_c111 bl_111 br_111 wl_105 vdd gnd cell_6t
Xbit_r106_c111 bl_111 br_111 wl_106 vdd gnd cell_6t
Xbit_r107_c111 bl_111 br_111 wl_107 vdd gnd cell_6t
Xbit_r108_c111 bl_111 br_111 wl_108 vdd gnd cell_6t
Xbit_r109_c111 bl_111 br_111 wl_109 vdd gnd cell_6t
Xbit_r110_c111 bl_111 br_111 wl_110 vdd gnd cell_6t
Xbit_r111_c111 bl_111 br_111 wl_111 vdd gnd cell_6t
Xbit_r112_c111 bl_111 br_111 wl_112 vdd gnd cell_6t
Xbit_r113_c111 bl_111 br_111 wl_113 vdd gnd cell_6t
Xbit_r114_c111 bl_111 br_111 wl_114 vdd gnd cell_6t
Xbit_r115_c111 bl_111 br_111 wl_115 vdd gnd cell_6t
Xbit_r116_c111 bl_111 br_111 wl_116 vdd gnd cell_6t
Xbit_r117_c111 bl_111 br_111 wl_117 vdd gnd cell_6t
Xbit_r118_c111 bl_111 br_111 wl_118 vdd gnd cell_6t
Xbit_r119_c111 bl_111 br_111 wl_119 vdd gnd cell_6t
Xbit_r120_c111 bl_111 br_111 wl_120 vdd gnd cell_6t
Xbit_r121_c111 bl_111 br_111 wl_121 vdd gnd cell_6t
Xbit_r122_c111 bl_111 br_111 wl_122 vdd gnd cell_6t
Xbit_r123_c111 bl_111 br_111 wl_123 vdd gnd cell_6t
Xbit_r124_c111 bl_111 br_111 wl_124 vdd gnd cell_6t
Xbit_r125_c111 bl_111 br_111 wl_125 vdd gnd cell_6t
Xbit_r126_c111 bl_111 br_111 wl_126 vdd gnd cell_6t
Xbit_r127_c111 bl_111 br_111 wl_127 vdd gnd cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd cell_6t
Xbit_r1_c112 bl_112 br_112 wl_1 vdd gnd cell_6t
Xbit_r2_c112 bl_112 br_112 wl_2 vdd gnd cell_6t
Xbit_r3_c112 bl_112 br_112 wl_3 vdd gnd cell_6t
Xbit_r4_c112 bl_112 br_112 wl_4 vdd gnd cell_6t
Xbit_r5_c112 bl_112 br_112 wl_5 vdd gnd cell_6t
Xbit_r6_c112 bl_112 br_112 wl_6 vdd gnd cell_6t
Xbit_r7_c112 bl_112 br_112 wl_7 vdd gnd cell_6t
Xbit_r8_c112 bl_112 br_112 wl_8 vdd gnd cell_6t
Xbit_r9_c112 bl_112 br_112 wl_9 vdd gnd cell_6t
Xbit_r10_c112 bl_112 br_112 wl_10 vdd gnd cell_6t
Xbit_r11_c112 bl_112 br_112 wl_11 vdd gnd cell_6t
Xbit_r12_c112 bl_112 br_112 wl_12 vdd gnd cell_6t
Xbit_r13_c112 bl_112 br_112 wl_13 vdd gnd cell_6t
Xbit_r14_c112 bl_112 br_112 wl_14 vdd gnd cell_6t
Xbit_r15_c112 bl_112 br_112 wl_15 vdd gnd cell_6t
Xbit_r16_c112 bl_112 br_112 wl_16 vdd gnd cell_6t
Xbit_r17_c112 bl_112 br_112 wl_17 vdd gnd cell_6t
Xbit_r18_c112 bl_112 br_112 wl_18 vdd gnd cell_6t
Xbit_r19_c112 bl_112 br_112 wl_19 vdd gnd cell_6t
Xbit_r20_c112 bl_112 br_112 wl_20 vdd gnd cell_6t
Xbit_r21_c112 bl_112 br_112 wl_21 vdd gnd cell_6t
Xbit_r22_c112 bl_112 br_112 wl_22 vdd gnd cell_6t
Xbit_r23_c112 bl_112 br_112 wl_23 vdd gnd cell_6t
Xbit_r24_c112 bl_112 br_112 wl_24 vdd gnd cell_6t
Xbit_r25_c112 bl_112 br_112 wl_25 vdd gnd cell_6t
Xbit_r26_c112 bl_112 br_112 wl_26 vdd gnd cell_6t
Xbit_r27_c112 bl_112 br_112 wl_27 vdd gnd cell_6t
Xbit_r28_c112 bl_112 br_112 wl_28 vdd gnd cell_6t
Xbit_r29_c112 bl_112 br_112 wl_29 vdd gnd cell_6t
Xbit_r30_c112 bl_112 br_112 wl_30 vdd gnd cell_6t
Xbit_r31_c112 bl_112 br_112 wl_31 vdd gnd cell_6t
Xbit_r32_c112 bl_112 br_112 wl_32 vdd gnd cell_6t
Xbit_r33_c112 bl_112 br_112 wl_33 vdd gnd cell_6t
Xbit_r34_c112 bl_112 br_112 wl_34 vdd gnd cell_6t
Xbit_r35_c112 bl_112 br_112 wl_35 vdd gnd cell_6t
Xbit_r36_c112 bl_112 br_112 wl_36 vdd gnd cell_6t
Xbit_r37_c112 bl_112 br_112 wl_37 vdd gnd cell_6t
Xbit_r38_c112 bl_112 br_112 wl_38 vdd gnd cell_6t
Xbit_r39_c112 bl_112 br_112 wl_39 vdd gnd cell_6t
Xbit_r40_c112 bl_112 br_112 wl_40 vdd gnd cell_6t
Xbit_r41_c112 bl_112 br_112 wl_41 vdd gnd cell_6t
Xbit_r42_c112 bl_112 br_112 wl_42 vdd gnd cell_6t
Xbit_r43_c112 bl_112 br_112 wl_43 vdd gnd cell_6t
Xbit_r44_c112 bl_112 br_112 wl_44 vdd gnd cell_6t
Xbit_r45_c112 bl_112 br_112 wl_45 vdd gnd cell_6t
Xbit_r46_c112 bl_112 br_112 wl_46 vdd gnd cell_6t
Xbit_r47_c112 bl_112 br_112 wl_47 vdd gnd cell_6t
Xbit_r48_c112 bl_112 br_112 wl_48 vdd gnd cell_6t
Xbit_r49_c112 bl_112 br_112 wl_49 vdd gnd cell_6t
Xbit_r50_c112 bl_112 br_112 wl_50 vdd gnd cell_6t
Xbit_r51_c112 bl_112 br_112 wl_51 vdd gnd cell_6t
Xbit_r52_c112 bl_112 br_112 wl_52 vdd gnd cell_6t
Xbit_r53_c112 bl_112 br_112 wl_53 vdd gnd cell_6t
Xbit_r54_c112 bl_112 br_112 wl_54 vdd gnd cell_6t
Xbit_r55_c112 bl_112 br_112 wl_55 vdd gnd cell_6t
Xbit_r56_c112 bl_112 br_112 wl_56 vdd gnd cell_6t
Xbit_r57_c112 bl_112 br_112 wl_57 vdd gnd cell_6t
Xbit_r58_c112 bl_112 br_112 wl_58 vdd gnd cell_6t
Xbit_r59_c112 bl_112 br_112 wl_59 vdd gnd cell_6t
Xbit_r60_c112 bl_112 br_112 wl_60 vdd gnd cell_6t
Xbit_r61_c112 bl_112 br_112 wl_61 vdd gnd cell_6t
Xbit_r62_c112 bl_112 br_112 wl_62 vdd gnd cell_6t
Xbit_r63_c112 bl_112 br_112 wl_63 vdd gnd cell_6t
Xbit_r64_c112 bl_112 br_112 wl_64 vdd gnd cell_6t
Xbit_r65_c112 bl_112 br_112 wl_65 vdd gnd cell_6t
Xbit_r66_c112 bl_112 br_112 wl_66 vdd gnd cell_6t
Xbit_r67_c112 bl_112 br_112 wl_67 vdd gnd cell_6t
Xbit_r68_c112 bl_112 br_112 wl_68 vdd gnd cell_6t
Xbit_r69_c112 bl_112 br_112 wl_69 vdd gnd cell_6t
Xbit_r70_c112 bl_112 br_112 wl_70 vdd gnd cell_6t
Xbit_r71_c112 bl_112 br_112 wl_71 vdd gnd cell_6t
Xbit_r72_c112 bl_112 br_112 wl_72 vdd gnd cell_6t
Xbit_r73_c112 bl_112 br_112 wl_73 vdd gnd cell_6t
Xbit_r74_c112 bl_112 br_112 wl_74 vdd gnd cell_6t
Xbit_r75_c112 bl_112 br_112 wl_75 vdd gnd cell_6t
Xbit_r76_c112 bl_112 br_112 wl_76 vdd gnd cell_6t
Xbit_r77_c112 bl_112 br_112 wl_77 vdd gnd cell_6t
Xbit_r78_c112 bl_112 br_112 wl_78 vdd gnd cell_6t
Xbit_r79_c112 bl_112 br_112 wl_79 vdd gnd cell_6t
Xbit_r80_c112 bl_112 br_112 wl_80 vdd gnd cell_6t
Xbit_r81_c112 bl_112 br_112 wl_81 vdd gnd cell_6t
Xbit_r82_c112 bl_112 br_112 wl_82 vdd gnd cell_6t
Xbit_r83_c112 bl_112 br_112 wl_83 vdd gnd cell_6t
Xbit_r84_c112 bl_112 br_112 wl_84 vdd gnd cell_6t
Xbit_r85_c112 bl_112 br_112 wl_85 vdd gnd cell_6t
Xbit_r86_c112 bl_112 br_112 wl_86 vdd gnd cell_6t
Xbit_r87_c112 bl_112 br_112 wl_87 vdd gnd cell_6t
Xbit_r88_c112 bl_112 br_112 wl_88 vdd gnd cell_6t
Xbit_r89_c112 bl_112 br_112 wl_89 vdd gnd cell_6t
Xbit_r90_c112 bl_112 br_112 wl_90 vdd gnd cell_6t
Xbit_r91_c112 bl_112 br_112 wl_91 vdd gnd cell_6t
Xbit_r92_c112 bl_112 br_112 wl_92 vdd gnd cell_6t
Xbit_r93_c112 bl_112 br_112 wl_93 vdd gnd cell_6t
Xbit_r94_c112 bl_112 br_112 wl_94 vdd gnd cell_6t
Xbit_r95_c112 bl_112 br_112 wl_95 vdd gnd cell_6t
Xbit_r96_c112 bl_112 br_112 wl_96 vdd gnd cell_6t
Xbit_r97_c112 bl_112 br_112 wl_97 vdd gnd cell_6t
Xbit_r98_c112 bl_112 br_112 wl_98 vdd gnd cell_6t
Xbit_r99_c112 bl_112 br_112 wl_99 vdd gnd cell_6t
Xbit_r100_c112 bl_112 br_112 wl_100 vdd gnd cell_6t
Xbit_r101_c112 bl_112 br_112 wl_101 vdd gnd cell_6t
Xbit_r102_c112 bl_112 br_112 wl_102 vdd gnd cell_6t
Xbit_r103_c112 bl_112 br_112 wl_103 vdd gnd cell_6t
Xbit_r104_c112 bl_112 br_112 wl_104 vdd gnd cell_6t
Xbit_r105_c112 bl_112 br_112 wl_105 vdd gnd cell_6t
Xbit_r106_c112 bl_112 br_112 wl_106 vdd gnd cell_6t
Xbit_r107_c112 bl_112 br_112 wl_107 vdd gnd cell_6t
Xbit_r108_c112 bl_112 br_112 wl_108 vdd gnd cell_6t
Xbit_r109_c112 bl_112 br_112 wl_109 vdd gnd cell_6t
Xbit_r110_c112 bl_112 br_112 wl_110 vdd gnd cell_6t
Xbit_r111_c112 bl_112 br_112 wl_111 vdd gnd cell_6t
Xbit_r112_c112 bl_112 br_112 wl_112 vdd gnd cell_6t
Xbit_r113_c112 bl_112 br_112 wl_113 vdd gnd cell_6t
Xbit_r114_c112 bl_112 br_112 wl_114 vdd gnd cell_6t
Xbit_r115_c112 bl_112 br_112 wl_115 vdd gnd cell_6t
Xbit_r116_c112 bl_112 br_112 wl_116 vdd gnd cell_6t
Xbit_r117_c112 bl_112 br_112 wl_117 vdd gnd cell_6t
Xbit_r118_c112 bl_112 br_112 wl_118 vdd gnd cell_6t
Xbit_r119_c112 bl_112 br_112 wl_119 vdd gnd cell_6t
Xbit_r120_c112 bl_112 br_112 wl_120 vdd gnd cell_6t
Xbit_r121_c112 bl_112 br_112 wl_121 vdd gnd cell_6t
Xbit_r122_c112 bl_112 br_112 wl_122 vdd gnd cell_6t
Xbit_r123_c112 bl_112 br_112 wl_123 vdd gnd cell_6t
Xbit_r124_c112 bl_112 br_112 wl_124 vdd gnd cell_6t
Xbit_r125_c112 bl_112 br_112 wl_125 vdd gnd cell_6t
Xbit_r126_c112 bl_112 br_112 wl_126 vdd gnd cell_6t
Xbit_r127_c112 bl_112 br_112 wl_127 vdd gnd cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd cell_6t
Xbit_r1_c113 bl_113 br_113 wl_1 vdd gnd cell_6t
Xbit_r2_c113 bl_113 br_113 wl_2 vdd gnd cell_6t
Xbit_r3_c113 bl_113 br_113 wl_3 vdd gnd cell_6t
Xbit_r4_c113 bl_113 br_113 wl_4 vdd gnd cell_6t
Xbit_r5_c113 bl_113 br_113 wl_5 vdd gnd cell_6t
Xbit_r6_c113 bl_113 br_113 wl_6 vdd gnd cell_6t
Xbit_r7_c113 bl_113 br_113 wl_7 vdd gnd cell_6t
Xbit_r8_c113 bl_113 br_113 wl_8 vdd gnd cell_6t
Xbit_r9_c113 bl_113 br_113 wl_9 vdd gnd cell_6t
Xbit_r10_c113 bl_113 br_113 wl_10 vdd gnd cell_6t
Xbit_r11_c113 bl_113 br_113 wl_11 vdd gnd cell_6t
Xbit_r12_c113 bl_113 br_113 wl_12 vdd gnd cell_6t
Xbit_r13_c113 bl_113 br_113 wl_13 vdd gnd cell_6t
Xbit_r14_c113 bl_113 br_113 wl_14 vdd gnd cell_6t
Xbit_r15_c113 bl_113 br_113 wl_15 vdd gnd cell_6t
Xbit_r16_c113 bl_113 br_113 wl_16 vdd gnd cell_6t
Xbit_r17_c113 bl_113 br_113 wl_17 vdd gnd cell_6t
Xbit_r18_c113 bl_113 br_113 wl_18 vdd gnd cell_6t
Xbit_r19_c113 bl_113 br_113 wl_19 vdd gnd cell_6t
Xbit_r20_c113 bl_113 br_113 wl_20 vdd gnd cell_6t
Xbit_r21_c113 bl_113 br_113 wl_21 vdd gnd cell_6t
Xbit_r22_c113 bl_113 br_113 wl_22 vdd gnd cell_6t
Xbit_r23_c113 bl_113 br_113 wl_23 vdd gnd cell_6t
Xbit_r24_c113 bl_113 br_113 wl_24 vdd gnd cell_6t
Xbit_r25_c113 bl_113 br_113 wl_25 vdd gnd cell_6t
Xbit_r26_c113 bl_113 br_113 wl_26 vdd gnd cell_6t
Xbit_r27_c113 bl_113 br_113 wl_27 vdd gnd cell_6t
Xbit_r28_c113 bl_113 br_113 wl_28 vdd gnd cell_6t
Xbit_r29_c113 bl_113 br_113 wl_29 vdd gnd cell_6t
Xbit_r30_c113 bl_113 br_113 wl_30 vdd gnd cell_6t
Xbit_r31_c113 bl_113 br_113 wl_31 vdd gnd cell_6t
Xbit_r32_c113 bl_113 br_113 wl_32 vdd gnd cell_6t
Xbit_r33_c113 bl_113 br_113 wl_33 vdd gnd cell_6t
Xbit_r34_c113 bl_113 br_113 wl_34 vdd gnd cell_6t
Xbit_r35_c113 bl_113 br_113 wl_35 vdd gnd cell_6t
Xbit_r36_c113 bl_113 br_113 wl_36 vdd gnd cell_6t
Xbit_r37_c113 bl_113 br_113 wl_37 vdd gnd cell_6t
Xbit_r38_c113 bl_113 br_113 wl_38 vdd gnd cell_6t
Xbit_r39_c113 bl_113 br_113 wl_39 vdd gnd cell_6t
Xbit_r40_c113 bl_113 br_113 wl_40 vdd gnd cell_6t
Xbit_r41_c113 bl_113 br_113 wl_41 vdd gnd cell_6t
Xbit_r42_c113 bl_113 br_113 wl_42 vdd gnd cell_6t
Xbit_r43_c113 bl_113 br_113 wl_43 vdd gnd cell_6t
Xbit_r44_c113 bl_113 br_113 wl_44 vdd gnd cell_6t
Xbit_r45_c113 bl_113 br_113 wl_45 vdd gnd cell_6t
Xbit_r46_c113 bl_113 br_113 wl_46 vdd gnd cell_6t
Xbit_r47_c113 bl_113 br_113 wl_47 vdd gnd cell_6t
Xbit_r48_c113 bl_113 br_113 wl_48 vdd gnd cell_6t
Xbit_r49_c113 bl_113 br_113 wl_49 vdd gnd cell_6t
Xbit_r50_c113 bl_113 br_113 wl_50 vdd gnd cell_6t
Xbit_r51_c113 bl_113 br_113 wl_51 vdd gnd cell_6t
Xbit_r52_c113 bl_113 br_113 wl_52 vdd gnd cell_6t
Xbit_r53_c113 bl_113 br_113 wl_53 vdd gnd cell_6t
Xbit_r54_c113 bl_113 br_113 wl_54 vdd gnd cell_6t
Xbit_r55_c113 bl_113 br_113 wl_55 vdd gnd cell_6t
Xbit_r56_c113 bl_113 br_113 wl_56 vdd gnd cell_6t
Xbit_r57_c113 bl_113 br_113 wl_57 vdd gnd cell_6t
Xbit_r58_c113 bl_113 br_113 wl_58 vdd gnd cell_6t
Xbit_r59_c113 bl_113 br_113 wl_59 vdd gnd cell_6t
Xbit_r60_c113 bl_113 br_113 wl_60 vdd gnd cell_6t
Xbit_r61_c113 bl_113 br_113 wl_61 vdd gnd cell_6t
Xbit_r62_c113 bl_113 br_113 wl_62 vdd gnd cell_6t
Xbit_r63_c113 bl_113 br_113 wl_63 vdd gnd cell_6t
Xbit_r64_c113 bl_113 br_113 wl_64 vdd gnd cell_6t
Xbit_r65_c113 bl_113 br_113 wl_65 vdd gnd cell_6t
Xbit_r66_c113 bl_113 br_113 wl_66 vdd gnd cell_6t
Xbit_r67_c113 bl_113 br_113 wl_67 vdd gnd cell_6t
Xbit_r68_c113 bl_113 br_113 wl_68 vdd gnd cell_6t
Xbit_r69_c113 bl_113 br_113 wl_69 vdd gnd cell_6t
Xbit_r70_c113 bl_113 br_113 wl_70 vdd gnd cell_6t
Xbit_r71_c113 bl_113 br_113 wl_71 vdd gnd cell_6t
Xbit_r72_c113 bl_113 br_113 wl_72 vdd gnd cell_6t
Xbit_r73_c113 bl_113 br_113 wl_73 vdd gnd cell_6t
Xbit_r74_c113 bl_113 br_113 wl_74 vdd gnd cell_6t
Xbit_r75_c113 bl_113 br_113 wl_75 vdd gnd cell_6t
Xbit_r76_c113 bl_113 br_113 wl_76 vdd gnd cell_6t
Xbit_r77_c113 bl_113 br_113 wl_77 vdd gnd cell_6t
Xbit_r78_c113 bl_113 br_113 wl_78 vdd gnd cell_6t
Xbit_r79_c113 bl_113 br_113 wl_79 vdd gnd cell_6t
Xbit_r80_c113 bl_113 br_113 wl_80 vdd gnd cell_6t
Xbit_r81_c113 bl_113 br_113 wl_81 vdd gnd cell_6t
Xbit_r82_c113 bl_113 br_113 wl_82 vdd gnd cell_6t
Xbit_r83_c113 bl_113 br_113 wl_83 vdd gnd cell_6t
Xbit_r84_c113 bl_113 br_113 wl_84 vdd gnd cell_6t
Xbit_r85_c113 bl_113 br_113 wl_85 vdd gnd cell_6t
Xbit_r86_c113 bl_113 br_113 wl_86 vdd gnd cell_6t
Xbit_r87_c113 bl_113 br_113 wl_87 vdd gnd cell_6t
Xbit_r88_c113 bl_113 br_113 wl_88 vdd gnd cell_6t
Xbit_r89_c113 bl_113 br_113 wl_89 vdd gnd cell_6t
Xbit_r90_c113 bl_113 br_113 wl_90 vdd gnd cell_6t
Xbit_r91_c113 bl_113 br_113 wl_91 vdd gnd cell_6t
Xbit_r92_c113 bl_113 br_113 wl_92 vdd gnd cell_6t
Xbit_r93_c113 bl_113 br_113 wl_93 vdd gnd cell_6t
Xbit_r94_c113 bl_113 br_113 wl_94 vdd gnd cell_6t
Xbit_r95_c113 bl_113 br_113 wl_95 vdd gnd cell_6t
Xbit_r96_c113 bl_113 br_113 wl_96 vdd gnd cell_6t
Xbit_r97_c113 bl_113 br_113 wl_97 vdd gnd cell_6t
Xbit_r98_c113 bl_113 br_113 wl_98 vdd gnd cell_6t
Xbit_r99_c113 bl_113 br_113 wl_99 vdd gnd cell_6t
Xbit_r100_c113 bl_113 br_113 wl_100 vdd gnd cell_6t
Xbit_r101_c113 bl_113 br_113 wl_101 vdd gnd cell_6t
Xbit_r102_c113 bl_113 br_113 wl_102 vdd gnd cell_6t
Xbit_r103_c113 bl_113 br_113 wl_103 vdd gnd cell_6t
Xbit_r104_c113 bl_113 br_113 wl_104 vdd gnd cell_6t
Xbit_r105_c113 bl_113 br_113 wl_105 vdd gnd cell_6t
Xbit_r106_c113 bl_113 br_113 wl_106 vdd gnd cell_6t
Xbit_r107_c113 bl_113 br_113 wl_107 vdd gnd cell_6t
Xbit_r108_c113 bl_113 br_113 wl_108 vdd gnd cell_6t
Xbit_r109_c113 bl_113 br_113 wl_109 vdd gnd cell_6t
Xbit_r110_c113 bl_113 br_113 wl_110 vdd gnd cell_6t
Xbit_r111_c113 bl_113 br_113 wl_111 vdd gnd cell_6t
Xbit_r112_c113 bl_113 br_113 wl_112 vdd gnd cell_6t
Xbit_r113_c113 bl_113 br_113 wl_113 vdd gnd cell_6t
Xbit_r114_c113 bl_113 br_113 wl_114 vdd gnd cell_6t
Xbit_r115_c113 bl_113 br_113 wl_115 vdd gnd cell_6t
Xbit_r116_c113 bl_113 br_113 wl_116 vdd gnd cell_6t
Xbit_r117_c113 bl_113 br_113 wl_117 vdd gnd cell_6t
Xbit_r118_c113 bl_113 br_113 wl_118 vdd gnd cell_6t
Xbit_r119_c113 bl_113 br_113 wl_119 vdd gnd cell_6t
Xbit_r120_c113 bl_113 br_113 wl_120 vdd gnd cell_6t
Xbit_r121_c113 bl_113 br_113 wl_121 vdd gnd cell_6t
Xbit_r122_c113 bl_113 br_113 wl_122 vdd gnd cell_6t
Xbit_r123_c113 bl_113 br_113 wl_123 vdd gnd cell_6t
Xbit_r124_c113 bl_113 br_113 wl_124 vdd gnd cell_6t
Xbit_r125_c113 bl_113 br_113 wl_125 vdd gnd cell_6t
Xbit_r126_c113 bl_113 br_113 wl_126 vdd gnd cell_6t
Xbit_r127_c113 bl_113 br_113 wl_127 vdd gnd cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd cell_6t
Xbit_r1_c114 bl_114 br_114 wl_1 vdd gnd cell_6t
Xbit_r2_c114 bl_114 br_114 wl_2 vdd gnd cell_6t
Xbit_r3_c114 bl_114 br_114 wl_3 vdd gnd cell_6t
Xbit_r4_c114 bl_114 br_114 wl_4 vdd gnd cell_6t
Xbit_r5_c114 bl_114 br_114 wl_5 vdd gnd cell_6t
Xbit_r6_c114 bl_114 br_114 wl_6 vdd gnd cell_6t
Xbit_r7_c114 bl_114 br_114 wl_7 vdd gnd cell_6t
Xbit_r8_c114 bl_114 br_114 wl_8 vdd gnd cell_6t
Xbit_r9_c114 bl_114 br_114 wl_9 vdd gnd cell_6t
Xbit_r10_c114 bl_114 br_114 wl_10 vdd gnd cell_6t
Xbit_r11_c114 bl_114 br_114 wl_11 vdd gnd cell_6t
Xbit_r12_c114 bl_114 br_114 wl_12 vdd gnd cell_6t
Xbit_r13_c114 bl_114 br_114 wl_13 vdd gnd cell_6t
Xbit_r14_c114 bl_114 br_114 wl_14 vdd gnd cell_6t
Xbit_r15_c114 bl_114 br_114 wl_15 vdd gnd cell_6t
Xbit_r16_c114 bl_114 br_114 wl_16 vdd gnd cell_6t
Xbit_r17_c114 bl_114 br_114 wl_17 vdd gnd cell_6t
Xbit_r18_c114 bl_114 br_114 wl_18 vdd gnd cell_6t
Xbit_r19_c114 bl_114 br_114 wl_19 vdd gnd cell_6t
Xbit_r20_c114 bl_114 br_114 wl_20 vdd gnd cell_6t
Xbit_r21_c114 bl_114 br_114 wl_21 vdd gnd cell_6t
Xbit_r22_c114 bl_114 br_114 wl_22 vdd gnd cell_6t
Xbit_r23_c114 bl_114 br_114 wl_23 vdd gnd cell_6t
Xbit_r24_c114 bl_114 br_114 wl_24 vdd gnd cell_6t
Xbit_r25_c114 bl_114 br_114 wl_25 vdd gnd cell_6t
Xbit_r26_c114 bl_114 br_114 wl_26 vdd gnd cell_6t
Xbit_r27_c114 bl_114 br_114 wl_27 vdd gnd cell_6t
Xbit_r28_c114 bl_114 br_114 wl_28 vdd gnd cell_6t
Xbit_r29_c114 bl_114 br_114 wl_29 vdd gnd cell_6t
Xbit_r30_c114 bl_114 br_114 wl_30 vdd gnd cell_6t
Xbit_r31_c114 bl_114 br_114 wl_31 vdd gnd cell_6t
Xbit_r32_c114 bl_114 br_114 wl_32 vdd gnd cell_6t
Xbit_r33_c114 bl_114 br_114 wl_33 vdd gnd cell_6t
Xbit_r34_c114 bl_114 br_114 wl_34 vdd gnd cell_6t
Xbit_r35_c114 bl_114 br_114 wl_35 vdd gnd cell_6t
Xbit_r36_c114 bl_114 br_114 wl_36 vdd gnd cell_6t
Xbit_r37_c114 bl_114 br_114 wl_37 vdd gnd cell_6t
Xbit_r38_c114 bl_114 br_114 wl_38 vdd gnd cell_6t
Xbit_r39_c114 bl_114 br_114 wl_39 vdd gnd cell_6t
Xbit_r40_c114 bl_114 br_114 wl_40 vdd gnd cell_6t
Xbit_r41_c114 bl_114 br_114 wl_41 vdd gnd cell_6t
Xbit_r42_c114 bl_114 br_114 wl_42 vdd gnd cell_6t
Xbit_r43_c114 bl_114 br_114 wl_43 vdd gnd cell_6t
Xbit_r44_c114 bl_114 br_114 wl_44 vdd gnd cell_6t
Xbit_r45_c114 bl_114 br_114 wl_45 vdd gnd cell_6t
Xbit_r46_c114 bl_114 br_114 wl_46 vdd gnd cell_6t
Xbit_r47_c114 bl_114 br_114 wl_47 vdd gnd cell_6t
Xbit_r48_c114 bl_114 br_114 wl_48 vdd gnd cell_6t
Xbit_r49_c114 bl_114 br_114 wl_49 vdd gnd cell_6t
Xbit_r50_c114 bl_114 br_114 wl_50 vdd gnd cell_6t
Xbit_r51_c114 bl_114 br_114 wl_51 vdd gnd cell_6t
Xbit_r52_c114 bl_114 br_114 wl_52 vdd gnd cell_6t
Xbit_r53_c114 bl_114 br_114 wl_53 vdd gnd cell_6t
Xbit_r54_c114 bl_114 br_114 wl_54 vdd gnd cell_6t
Xbit_r55_c114 bl_114 br_114 wl_55 vdd gnd cell_6t
Xbit_r56_c114 bl_114 br_114 wl_56 vdd gnd cell_6t
Xbit_r57_c114 bl_114 br_114 wl_57 vdd gnd cell_6t
Xbit_r58_c114 bl_114 br_114 wl_58 vdd gnd cell_6t
Xbit_r59_c114 bl_114 br_114 wl_59 vdd gnd cell_6t
Xbit_r60_c114 bl_114 br_114 wl_60 vdd gnd cell_6t
Xbit_r61_c114 bl_114 br_114 wl_61 vdd gnd cell_6t
Xbit_r62_c114 bl_114 br_114 wl_62 vdd gnd cell_6t
Xbit_r63_c114 bl_114 br_114 wl_63 vdd gnd cell_6t
Xbit_r64_c114 bl_114 br_114 wl_64 vdd gnd cell_6t
Xbit_r65_c114 bl_114 br_114 wl_65 vdd gnd cell_6t
Xbit_r66_c114 bl_114 br_114 wl_66 vdd gnd cell_6t
Xbit_r67_c114 bl_114 br_114 wl_67 vdd gnd cell_6t
Xbit_r68_c114 bl_114 br_114 wl_68 vdd gnd cell_6t
Xbit_r69_c114 bl_114 br_114 wl_69 vdd gnd cell_6t
Xbit_r70_c114 bl_114 br_114 wl_70 vdd gnd cell_6t
Xbit_r71_c114 bl_114 br_114 wl_71 vdd gnd cell_6t
Xbit_r72_c114 bl_114 br_114 wl_72 vdd gnd cell_6t
Xbit_r73_c114 bl_114 br_114 wl_73 vdd gnd cell_6t
Xbit_r74_c114 bl_114 br_114 wl_74 vdd gnd cell_6t
Xbit_r75_c114 bl_114 br_114 wl_75 vdd gnd cell_6t
Xbit_r76_c114 bl_114 br_114 wl_76 vdd gnd cell_6t
Xbit_r77_c114 bl_114 br_114 wl_77 vdd gnd cell_6t
Xbit_r78_c114 bl_114 br_114 wl_78 vdd gnd cell_6t
Xbit_r79_c114 bl_114 br_114 wl_79 vdd gnd cell_6t
Xbit_r80_c114 bl_114 br_114 wl_80 vdd gnd cell_6t
Xbit_r81_c114 bl_114 br_114 wl_81 vdd gnd cell_6t
Xbit_r82_c114 bl_114 br_114 wl_82 vdd gnd cell_6t
Xbit_r83_c114 bl_114 br_114 wl_83 vdd gnd cell_6t
Xbit_r84_c114 bl_114 br_114 wl_84 vdd gnd cell_6t
Xbit_r85_c114 bl_114 br_114 wl_85 vdd gnd cell_6t
Xbit_r86_c114 bl_114 br_114 wl_86 vdd gnd cell_6t
Xbit_r87_c114 bl_114 br_114 wl_87 vdd gnd cell_6t
Xbit_r88_c114 bl_114 br_114 wl_88 vdd gnd cell_6t
Xbit_r89_c114 bl_114 br_114 wl_89 vdd gnd cell_6t
Xbit_r90_c114 bl_114 br_114 wl_90 vdd gnd cell_6t
Xbit_r91_c114 bl_114 br_114 wl_91 vdd gnd cell_6t
Xbit_r92_c114 bl_114 br_114 wl_92 vdd gnd cell_6t
Xbit_r93_c114 bl_114 br_114 wl_93 vdd gnd cell_6t
Xbit_r94_c114 bl_114 br_114 wl_94 vdd gnd cell_6t
Xbit_r95_c114 bl_114 br_114 wl_95 vdd gnd cell_6t
Xbit_r96_c114 bl_114 br_114 wl_96 vdd gnd cell_6t
Xbit_r97_c114 bl_114 br_114 wl_97 vdd gnd cell_6t
Xbit_r98_c114 bl_114 br_114 wl_98 vdd gnd cell_6t
Xbit_r99_c114 bl_114 br_114 wl_99 vdd gnd cell_6t
Xbit_r100_c114 bl_114 br_114 wl_100 vdd gnd cell_6t
Xbit_r101_c114 bl_114 br_114 wl_101 vdd gnd cell_6t
Xbit_r102_c114 bl_114 br_114 wl_102 vdd gnd cell_6t
Xbit_r103_c114 bl_114 br_114 wl_103 vdd gnd cell_6t
Xbit_r104_c114 bl_114 br_114 wl_104 vdd gnd cell_6t
Xbit_r105_c114 bl_114 br_114 wl_105 vdd gnd cell_6t
Xbit_r106_c114 bl_114 br_114 wl_106 vdd gnd cell_6t
Xbit_r107_c114 bl_114 br_114 wl_107 vdd gnd cell_6t
Xbit_r108_c114 bl_114 br_114 wl_108 vdd gnd cell_6t
Xbit_r109_c114 bl_114 br_114 wl_109 vdd gnd cell_6t
Xbit_r110_c114 bl_114 br_114 wl_110 vdd gnd cell_6t
Xbit_r111_c114 bl_114 br_114 wl_111 vdd gnd cell_6t
Xbit_r112_c114 bl_114 br_114 wl_112 vdd gnd cell_6t
Xbit_r113_c114 bl_114 br_114 wl_113 vdd gnd cell_6t
Xbit_r114_c114 bl_114 br_114 wl_114 vdd gnd cell_6t
Xbit_r115_c114 bl_114 br_114 wl_115 vdd gnd cell_6t
Xbit_r116_c114 bl_114 br_114 wl_116 vdd gnd cell_6t
Xbit_r117_c114 bl_114 br_114 wl_117 vdd gnd cell_6t
Xbit_r118_c114 bl_114 br_114 wl_118 vdd gnd cell_6t
Xbit_r119_c114 bl_114 br_114 wl_119 vdd gnd cell_6t
Xbit_r120_c114 bl_114 br_114 wl_120 vdd gnd cell_6t
Xbit_r121_c114 bl_114 br_114 wl_121 vdd gnd cell_6t
Xbit_r122_c114 bl_114 br_114 wl_122 vdd gnd cell_6t
Xbit_r123_c114 bl_114 br_114 wl_123 vdd gnd cell_6t
Xbit_r124_c114 bl_114 br_114 wl_124 vdd gnd cell_6t
Xbit_r125_c114 bl_114 br_114 wl_125 vdd gnd cell_6t
Xbit_r126_c114 bl_114 br_114 wl_126 vdd gnd cell_6t
Xbit_r127_c114 bl_114 br_114 wl_127 vdd gnd cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd cell_6t
Xbit_r1_c115 bl_115 br_115 wl_1 vdd gnd cell_6t
Xbit_r2_c115 bl_115 br_115 wl_2 vdd gnd cell_6t
Xbit_r3_c115 bl_115 br_115 wl_3 vdd gnd cell_6t
Xbit_r4_c115 bl_115 br_115 wl_4 vdd gnd cell_6t
Xbit_r5_c115 bl_115 br_115 wl_5 vdd gnd cell_6t
Xbit_r6_c115 bl_115 br_115 wl_6 vdd gnd cell_6t
Xbit_r7_c115 bl_115 br_115 wl_7 vdd gnd cell_6t
Xbit_r8_c115 bl_115 br_115 wl_8 vdd gnd cell_6t
Xbit_r9_c115 bl_115 br_115 wl_9 vdd gnd cell_6t
Xbit_r10_c115 bl_115 br_115 wl_10 vdd gnd cell_6t
Xbit_r11_c115 bl_115 br_115 wl_11 vdd gnd cell_6t
Xbit_r12_c115 bl_115 br_115 wl_12 vdd gnd cell_6t
Xbit_r13_c115 bl_115 br_115 wl_13 vdd gnd cell_6t
Xbit_r14_c115 bl_115 br_115 wl_14 vdd gnd cell_6t
Xbit_r15_c115 bl_115 br_115 wl_15 vdd gnd cell_6t
Xbit_r16_c115 bl_115 br_115 wl_16 vdd gnd cell_6t
Xbit_r17_c115 bl_115 br_115 wl_17 vdd gnd cell_6t
Xbit_r18_c115 bl_115 br_115 wl_18 vdd gnd cell_6t
Xbit_r19_c115 bl_115 br_115 wl_19 vdd gnd cell_6t
Xbit_r20_c115 bl_115 br_115 wl_20 vdd gnd cell_6t
Xbit_r21_c115 bl_115 br_115 wl_21 vdd gnd cell_6t
Xbit_r22_c115 bl_115 br_115 wl_22 vdd gnd cell_6t
Xbit_r23_c115 bl_115 br_115 wl_23 vdd gnd cell_6t
Xbit_r24_c115 bl_115 br_115 wl_24 vdd gnd cell_6t
Xbit_r25_c115 bl_115 br_115 wl_25 vdd gnd cell_6t
Xbit_r26_c115 bl_115 br_115 wl_26 vdd gnd cell_6t
Xbit_r27_c115 bl_115 br_115 wl_27 vdd gnd cell_6t
Xbit_r28_c115 bl_115 br_115 wl_28 vdd gnd cell_6t
Xbit_r29_c115 bl_115 br_115 wl_29 vdd gnd cell_6t
Xbit_r30_c115 bl_115 br_115 wl_30 vdd gnd cell_6t
Xbit_r31_c115 bl_115 br_115 wl_31 vdd gnd cell_6t
Xbit_r32_c115 bl_115 br_115 wl_32 vdd gnd cell_6t
Xbit_r33_c115 bl_115 br_115 wl_33 vdd gnd cell_6t
Xbit_r34_c115 bl_115 br_115 wl_34 vdd gnd cell_6t
Xbit_r35_c115 bl_115 br_115 wl_35 vdd gnd cell_6t
Xbit_r36_c115 bl_115 br_115 wl_36 vdd gnd cell_6t
Xbit_r37_c115 bl_115 br_115 wl_37 vdd gnd cell_6t
Xbit_r38_c115 bl_115 br_115 wl_38 vdd gnd cell_6t
Xbit_r39_c115 bl_115 br_115 wl_39 vdd gnd cell_6t
Xbit_r40_c115 bl_115 br_115 wl_40 vdd gnd cell_6t
Xbit_r41_c115 bl_115 br_115 wl_41 vdd gnd cell_6t
Xbit_r42_c115 bl_115 br_115 wl_42 vdd gnd cell_6t
Xbit_r43_c115 bl_115 br_115 wl_43 vdd gnd cell_6t
Xbit_r44_c115 bl_115 br_115 wl_44 vdd gnd cell_6t
Xbit_r45_c115 bl_115 br_115 wl_45 vdd gnd cell_6t
Xbit_r46_c115 bl_115 br_115 wl_46 vdd gnd cell_6t
Xbit_r47_c115 bl_115 br_115 wl_47 vdd gnd cell_6t
Xbit_r48_c115 bl_115 br_115 wl_48 vdd gnd cell_6t
Xbit_r49_c115 bl_115 br_115 wl_49 vdd gnd cell_6t
Xbit_r50_c115 bl_115 br_115 wl_50 vdd gnd cell_6t
Xbit_r51_c115 bl_115 br_115 wl_51 vdd gnd cell_6t
Xbit_r52_c115 bl_115 br_115 wl_52 vdd gnd cell_6t
Xbit_r53_c115 bl_115 br_115 wl_53 vdd gnd cell_6t
Xbit_r54_c115 bl_115 br_115 wl_54 vdd gnd cell_6t
Xbit_r55_c115 bl_115 br_115 wl_55 vdd gnd cell_6t
Xbit_r56_c115 bl_115 br_115 wl_56 vdd gnd cell_6t
Xbit_r57_c115 bl_115 br_115 wl_57 vdd gnd cell_6t
Xbit_r58_c115 bl_115 br_115 wl_58 vdd gnd cell_6t
Xbit_r59_c115 bl_115 br_115 wl_59 vdd gnd cell_6t
Xbit_r60_c115 bl_115 br_115 wl_60 vdd gnd cell_6t
Xbit_r61_c115 bl_115 br_115 wl_61 vdd gnd cell_6t
Xbit_r62_c115 bl_115 br_115 wl_62 vdd gnd cell_6t
Xbit_r63_c115 bl_115 br_115 wl_63 vdd gnd cell_6t
Xbit_r64_c115 bl_115 br_115 wl_64 vdd gnd cell_6t
Xbit_r65_c115 bl_115 br_115 wl_65 vdd gnd cell_6t
Xbit_r66_c115 bl_115 br_115 wl_66 vdd gnd cell_6t
Xbit_r67_c115 bl_115 br_115 wl_67 vdd gnd cell_6t
Xbit_r68_c115 bl_115 br_115 wl_68 vdd gnd cell_6t
Xbit_r69_c115 bl_115 br_115 wl_69 vdd gnd cell_6t
Xbit_r70_c115 bl_115 br_115 wl_70 vdd gnd cell_6t
Xbit_r71_c115 bl_115 br_115 wl_71 vdd gnd cell_6t
Xbit_r72_c115 bl_115 br_115 wl_72 vdd gnd cell_6t
Xbit_r73_c115 bl_115 br_115 wl_73 vdd gnd cell_6t
Xbit_r74_c115 bl_115 br_115 wl_74 vdd gnd cell_6t
Xbit_r75_c115 bl_115 br_115 wl_75 vdd gnd cell_6t
Xbit_r76_c115 bl_115 br_115 wl_76 vdd gnd cell_6t
Xbit_r77_c115 bl_115 br_115 wl_77 vdd gnd cell_6t
Xbit_r78_c115 bl_115 br_115 wl_78 vdd gnd cell_6t
Xbit_r79_c115 bl_115 br_115 wl_79 vdd gnd cell_6t
Xbit_r80_c115 bl_115 br_115 wl_80 vdd gnd cell_6t
Xbit_r81_c115 bl_115 br_115 wl_81 vdd gnd cell_6t
Xbit_r82_c115 bl_115 br_115 wl_82 vdd gnd cell_6t
Xbit_r83_c115 bl_115 br_115 wl_83 vdd gnd cell_6t
Xbit_r84_c115 bl_115 br_115 wl_84 vdd gnd cell_6t
Xbit_r85_c115 bl_115 br_115 wl_85 vdd gnd cell_6t
Xbit_r86_c115 bl_115 br_115 wl_86 vdd gnd cell_6t
Xbit_r87_c115 bl_115 br_115 wl_87 vdd gnd cell_6t
Xbit_r88_c115 bl_115 br_115 wl_88 vdd gnd cell_6t
Xbit_r89_c115 bl_115 br_115 wl_89 vdd gnd cell_6t
Xbit_r90_c115 bl_115 br_115 wl_90 vdd gnd cell_6t
Xbit_r91_c115 bl_115 br_115 wl_91 vdd gnd cell_6t
Xbit_r92_c115 bl_115 br_115 wl_92 vdd gnd cell_6t
Xbit_r93_c115 bl_115 br_115 wl_93 vdd gnd cell_6t
Xbit_r94_c115 bl_115 br_115 wl_94 vdd gnd cell_6t
Xbit_r95_c115 bl_115 br_115 wl_95 vdd gnd cell_6t
Xbit_r96_c115 bl_115 br_115 wl_96 vdd gnd cell_6t
Xbit_r97_c115 bl_115 br_115 wl_97 vdd gnd cell_6t
Xbit_r98_c115 bl_115 br_115 wl_98 vdd gnd cell_6t
Xbit_r99_c115 bl_115 br_115 wl_99 vdd gnd cell_6t
Xbit_r100_c115 bl_115 br_115 wl_100 vdd gnd cell_6t
Xbit_r101_c115 bl_115 br_115 wl_101 vdd gnd cell_6t
Xbit_r102_c115 bl_115 br_115 wl_102 vdd gnd cell_6t
Xbit_r103_c115 bl_115 br_115 wl_103 vdd gnd cell_6t
Xbit_r104_c115 bl_115 br_115 wl_104 vdd gnd cell_6t
Xbit_r105_c115 bl_115 br_115 wl_105 vdd gnd cell_6t
Xbit_r106_c115 bl_115 br_115 wl_106 vdd gnd cell_6t
Xbit_r107_c115 bl_115 br_115 wl_107 vdd gnd cell_6t
Xbit_r108_c115 bl_115 br_115 wl_108 vdd gnd cell_6t
Xbit_r109_c115 bl_115 br_115 wl_109 vdd gnd cell_6t
Xbit_r110_c115 bl_115 br_115 wl_110 vdd gnd cell_6t
Xbit_r111_c115 bl_115 br_115 wl_111 vdd gnd cell_6t
Xbit_r112_c115 bl_115 br_115 wl_112 vdd gnd cell_6t
Xbit_r113_c115 bl_115 br_115 wl_113 vdd gnd cell_6t
Xbit_r114_c115 bl_115 br_115 wl_114 vdd gnd cell_6t
Xbit_r115_c115 bl_115 br_115 wl_115 vdd gnd cell_6t
Xbit_r116_c115 bl_115 br_115 wl_116 vdd gnd cell_6t
Xbit_r117_c115 bl_115 br_115 wl_117 vdd gnd cell_6t
Xbit_r118_c115 bl_115 br_115 wl_118 vdd gnd cell_6t
Xbit_r119_c115 bl_115 br_115 wl_119 vdd gnd cell_6t
Xbit_r120_c115 bl_115 br_115 wl_120 vdd gnd cell_6t
Xbit_r121_c115 bl_115 br_115 wl_121 vdd gnd cell_6t
Xbit_r122_c115 bl_115 br_115 wl_122 vdd gnd cell_6t
Xbit_r123_c115 bl_115 br_115 wl_123 vdd gnd cell_6t
Xbit_r124_c115 bl_115 br_115 wl_124 vdd gnd cell_6t
Xbit_r125_c115 bl_115 br_115 wl_125 vdd gnd cell_6t
Xbit_r126_c115 bl_115 br_115 wl_126 vdd gnd cell_6t
Xbit_r127_c115 bl_115 br_115 wl_127 vdd gnd cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd cell_6t
Xbit_r1_c116 bl_116 br_116 wl_1 vdd gnd cell_6t
Xbit_r2_c116 bl_116 br_116 wl_2 vdd gnd cell_6t
Xbit_r3_c116 bl_116 br_116 wl_3 vdd gnd cell_6t
Xbit_r4_c116 bl_116 br_116 wl_4 vdd gnd cell_6t
Xbit_r5_c116 bl_116 br_116 wl_5 vdd gnd cell_6t
Xbit_r6_c116 bl_116 br_116 wl_6 vdd gnd cell_6t
Xbit_r7_c116 bl_116 br_116 wl_7 vdd gnd cell_6t
Xbit_r8_c116 bl_116 br_116 wl_8 vdd gnd cell_6t
Xbit_r9_c116 bl_116 br_116 wl_9 vdd gnd cell_6t
Xbit_r10_c116 bl_116 br_116 wl_10 vdd gnd cell_6t
Xbit_r11_c116 bl_116 br_116 wl_11 vdd gnd cell_6t
Xbit_r12_c116 bl_116 br_116 wl_12 vdd gnd cell_6t
Xbit_r13_c116 bl_116 br_116 wl_13 vdd gnd cell_6t
Xbit_r14_c116 bl_116 br_116 wl_14 vdd gnd cell_6t
Xbit_r15_c116 bl_116 br_116 wl_15 vdd gnd cell_6t
Xbit_r16_c116 bl_116 br_116 wl_16 vdd gnd cell_6t
Xbit_r17_c116 bl_116 br_116 wl_17 vdd gnd cell_6t
Xbit_r18_c116 bl_116 br_116 wl_18 vdd gnd cell_6t
Xbit_r19_c116 bl_116 br_116 wl_19 vdd gnd cell_6t
Xbit_r20_c116 bl_116 br_116 wl_20 vdd gnd cell_6t
Xbit_r21_c116 bl_116 br_116 wl_21 vdd gnd cell_6t
Xbit_r22_c116 bl_116 br_116 wl_22 vdd gnd cell_6t
Xbit_r23_c116 bl_116 br_116 wl_23 vdd gnd cell_6t
Xbit_r24_c116 bl_116 br_116 wl_24 vdd gnd cell_6t
Xbit_r25_c116 bl_116 br_116 wl_25 vdd gnd cell_6t
Xbit_r26_c116 bl_116 br_116 wl_26 vdd gnd cell_6t
Xbit_r27_c116 bl_116 br_116 wl_27 vdd gnd cell_6t
Xbit_r28_c116 bl_116 br_116 wl_28 vdd gnd cell_6t
Xbit_r29_c116 bl_116 br_116 wl_29 vdd gnd cell_6t
Xbit_r30_c116 bl_116 br_116 wl_30 vdd gnd cell_6t
Xbit_r31_c116 bl_116 br_116 wl_31 vdd gnd cell_6t
Xbit_r32_c116 bl_116 br_116 wl_32 vdd gnd cell_6t
Xbit_r33_c116 bl_116 br_116 wl_33 vdd gnd cell_6t
Xbit_r34_c116 bl_116 br_116 wl_34 vdd gnd cell_6t
Xbit_r35_c116 bl_116 br_116 wl_35 vdd gnd cell_6t
Xbit_r36_c116 bl_116 br_116 wl_36 vdd gnd cell_6t
Xbit_r37_c116 bl_116 br_116 wl_37 vdd gnd cell_6t
Xbit_r38_c116 bl_116 br_116 wl_38 vdd gnd cell_6t
Xbit_r39_c116 bl_116 br_116 wl_39 vdd gnd cell_6t
Xbit_r40_c116 bl_116 br_116 wl_40 vdd gnd cell_6t
Xbit_r41_c116 bl_116 br_116 wl_41 vdd gnd cell_6t
Xbit_r42_c116 bl_116 br_116 wl_42 vdd gnd cell_6t
Xbit_r43_c116 bl_116 br_116 wl_43 vdd gnd cell_6t
Xbit_r44_c116 bl_116 br_116 wl_44 vdd gnd cell_6t
Xbit_r45_c116 bl_116 br_116 wl_45 vdd gnd cell_6t
Xbit_r46_c116 bl_116 br_116 wl_46 vdd gnd cell_6t
Xbit_r47_c116 bl_116 br_116 wl_47 vdd gnd cell_6t
Xbit_r48_c116 bl_116 br_116 wl_48 vdd gnd cell_6t
Xbit_r49_c116 bl_116 br_116 wl_49 vdd gnd cell_6t
Xbit_r50_c116 bl_116 br_116 wl_50 vdd gnd cell_6t
Xbit_r51_c116 bl_116 br_116 wl_51 vdd gnd cell_6t
Xbit_r52_c116 bl_116 br_116 wl_52 vdd gnd cell_6t
Xbit_r53_c116 bl_116 br_116 wl_53 vdd gnd cell_6t
Xbit_r54_c116 bl_116 br_116 wl_54 vdd gnd cell_6t
Xbit_r55_c116 bl_116 br_116 wl_55 vdd gnd cell_6t
Xbit_r56_c116 bl_116 br_116 wl_56 vdd gnd cell_6t
Xbit_r57_c116 bl_116 br_116 wl_57 vdd gnd cell_6t
Xbit_r58_c116 bl_116 br_116 wl_58 vdd gnd cell_6t
Xbit_r59_c116 bl_116 br_116 wl_59 vdd gnd cell_6t
Xbit_r60_c116 bl_116 br_116 wl_60 vdd gnd cell_6t
Xbit_r61_c116 bl_116 br_116 wl_61 vdd gnd cell_6t
Xbit_r62_c116 bl_116 br_116 wl_62 vdd gnd cell_6t
Xbit_r63_c116 bl_116 br_116 wl_63 vdd gnd cell_6t
Xbit_r64_c116 bl_116 br_116 wl_64 vdd gnd cell_6t
Xbit_r65_c116 bl_116 br_116 wl_65 vdd gnd cell_6t
Xbit_r66_c116 bl_116 br_116 wl_66 vdd gnd cell_6t
Xbit_r67_c116 bl_116 br_116 wl_67 vdd gnd cell_6t
Xbit_r68_c116 bl_116 br_116 wl_68 vdd gnd cell_6t
Xbit_r69_c116 bl_116 br_116 wl_69 vdd gnd cell_6t
Xbit_r70_c116 bl_116 br_116 wl_70 vdd gnd cell_6t
Xbit_r71_c116 bl_116 br_116 wl_71 vdd gnd cell_6t
Xbit_r72_c116 bl_116 br_116 wl_72 vdd gnd cell_6t
Xbit_r73_c116 bl_116 br_116 wl_73 vdd gnd cell_6t
Xbit_r74_c116 bl_116 br_116 wl_74 vdd gnd cell_6t
Xbit_r75_c116 bl_116 br_116 wl_75 vdd gnd cell_6t
Xbit_r76_c116 bl_116 br_116 wl_76 vdd gnd cell_6t
Xbit_r77_c116 bl_116 br_116 wl_77 vdd gnd cell_6t
Xbit_r78_c116 bl_116 br_116 wl_78 vdd gnd cell_6t
Xbit_r79_c116 bl_116 br_116 wl_79 vdd gnd cell_6t
Xbit_r80_c116 bl_116 br_116 wl_80 vdd gnd cell_6t
Xbit_r81_c116 bl_116 br_116 wl_81 vdd gnd cell_6t
Xbit_r82_c116 bl_116 br_116 wl_82 vdd gnd cell_6t
Xbit_r83_c116 bl_116 br_116 wl_83 vdd gnd cell_6t
Xbit_r84_c116 bl_116 br_116 wl_84 vdd gnd cell_6t
Xbit_r85_c116 bl_116 br_116 wl_85 vdd gnd cell_6t
Xbit_r86_c116 bl_116 br_116 wl_86 vdd gnd cell_6t
Xbit_r87_c116 bl_116 br_116 wl_87 vdd gnd cell_6t
Xbit_r88_c116 bl_116 br_116 wl_88 vdd gnd cell_6t
Xbit_r89_c116 bl_116 br_116 wl_89 vdd gnd cell_6t
Xbit_r90_c116 bl_116 br_116 wl_90 vdd gnd cell_6t
Xbit_r91_c116 bl_116 br_116 wl_91 vdd gnd cell_6t
Xbit_r92_c116 bl_116 br_116 wl_92 vdd gnd cell_6t
Xbit_r93_c116 bl_116 br_116 wl_93 vdd gnd cell_6t
Xbit_r94_c116 bl_116 br_116 wl_94 vdd gnd cell_6t
Xbit_r95_c116 bl_116 br_116 wl_95 vdd gnd cell_6t
Xbit_r96_c116 bl_116 br_116 wl_96 vdd gnd cell_6t
Xbit_r97_c116 bl_116 br_116 wl_97 vdd gnd cell_6t
Xbit_r98_c116 bl_116 br_116 wl_98 vdd gnd cell_6t
Xbit_r99_c116 bl_116 br_116 wl_99 vdd gnd cell_6t
Xbit_r100_c116 bl_116 br_116 wl_100 vdd gnd cell_6t
Xbit_r101_c116 bl_116 br_116 wl_101 vdd gnd cell_6t
Xbit_r102_c116 bl_116 br_116 wl_102 vdd gnd cell_6t
Xbit_r103_c116 bl_116 br_116 wl_103 vdd gnd cell_6t
Xbit_r104_c116 bl_116 br_116 wl_104 vdd gnd cell_6t
Xbit_r105_c116 bl_116 br_116 wl_105 vdd gnd cell_6t
Xbit_r106_c116 bl_116 br_116 wl_106 vdd gnd cell_6t
Xbit_r107_c116 bl_116 br_116 wl_107 vdd gnd cell_6t
Xbit_r108_c116 bl_116 br_116 wl_108 vdd gnd cell_6t
Xbit_r109_c116 bl_116 br_116 wl_109 vdd gnd cell_6t
Xbit_r110_c116 bl_116 br_116 wl_110 vdd gnd cell_6t
Xbit_r111_c116 bl_116 br_116 wl_111 vdd gnd cell_6t
Xbit_r112_c116 bl_116 br_116 wl_112 vdd gnd cell_6t
Xbit_r113_c116 bl_116 br_116 wl_113 vdd gnd cell_6t
Xbit_r114_c116 bl_116 br_116 wl_114 vdd gnd cell_6t
Xbit_r115_c116 bl_116 br_116 wl_115 vdd gnd cell_6t
Xbit_r116_c116 bl_116 br_116 wl_116 vdd gnd cell_6t
Xbit_r117_c116 bl_116 br_116 wl_117 vdd gnd cell_6t
Xbit_r118_c116 bl_116 br_116 wl_118 vdd gnd cell_6t
Xbit_r119_c116 bl_116 br_116 wl_119 vdd gnd cell_6t
Xbit_r120_c116 bl_116 br_116 wl_120 vdd gnd cell_6t
Xbit_r121_c116 bl_116 br_116 wl_121 vdd gnd cell_6t
Xbit_r122_c116 bl_116 br_116 wl_122 vdd gnd cell_6t
Xbit_r123_c116 bl_116 br_116 wl_123 vdd gnd cell_6t
Xbit_r124_c116 bl_116 br_116 wl_124 vdd gnd cell_6t
Xbit_r125_c116 bl_116 br_116 wl_125 vdd gnd cell_6t
Xbit_r126_c116 bl_116 br_116 wl_126 vdd gnd cell_6t
Xbit_r127_c116 bl_116 br_116 wl_127 vdd gnd cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd cell_6t
Xbit_r1_c117 bl_117 br_117 wl_1 vdd gnd cell_6t
Xbit_r2_c117 bl_117 br_117 wl_2 vdd gnd cell_6t
Xbit_r3_c117 bl_117 br_117 wl_3 vdd gnd cell_6t
Xbit_r4_c117 bl_117 br_117 wl_4 vdd gnd cell_6t
Xbit_r5_c117 bl_117 br_117 wl_5 vdd gnd cell_6t
Xbit_r6_c117 bl_117 br_117 wl_6 vdd gnd cell_6t
Xbit_r7_c117 bl_117 br_117 wl_7 vdd gnd cell_6t
Xbit_r8_c117 bl_117 br_117 wl_8 vdd gnd cell_6t
Xbit_r9_c117 bl_117 br_117 wl_9 vdd gnd cell_6t
Xbit_r10_c117 bl_117 br_117 wl_10 vdd gnd cell_6t
Xbit_r11_c117 bl_117 br_117 wl_11 vdd gnd cell_6t
Xbit_r12_c117 bl_117 br_117 wl_12 vdd gnd cell_6t
Xbit_r13_c117 bl_117 br_117 wl_13 vdd gnd cell_6t
Xbit_r14_c117 bl_117 br_117 wl_14 vdd gnd cell_6t
Xbit_r15_c117 bl_117 br_117 wl_15 vdd gnd cell_6t
Xbit_r16_c117 bl_117 br_117 wl_16 vdd gnd cell_6t
Xbit_r17_c117 bl_117 br_117 wl_17 vdd gnd cell_6t
Xbit_r18_c117 bl_117 br_117 wl_18 vdd gnd cell_6t
Xbit_r19_c117 bl_117 br_117 wl_19 vdd gnd cell_6t
Xbit_r20_c117 bl_117 br_117 wl_20 vdd gnd cell_6t
Xbit_r21_c117 bl_117 br_117 wl_21 vdd gnd cell_6t
Xbit_r22_c117 bl_117 br_117 wl_22 vdd gnd cell_6t
Xbit_r23_c117 bl_117 br_117 wl_23 vdd gnd cell_6t
Xbit_r24_c117 bl_117 br_117 wl_24 vdd gnd cell_6t
Xbit_r25_c117 bl_117 br_117 wl_25 vdd gnd cell_6t
Xbit_r26_c117 bl_117 br_117 wl_26 vdd gnd cell_6t
Xbit_r27_c117 bl_117 br_117 wl_27 vdd gnd cell_6t
Xbit_r28_c117 bl_117 br_117 wl_28 vdd gnd cell_6t
Xbit_r29_c117 bl_117 br_117 wl_29 vdd gnd cell_6t
Xbit_r30_c117 bl_117 br_117 wl_30 vdd gnd cell_6t
Xbit_r31_c117 bl_117 br_117 wl_31 vdd gnd cell_6t
Xbit_r32_c117 bl_117 br_117 wl_32 vdd gnd cell_6t
Xbit_r33_c117 bl_117 br_117 wl_33 vdd gnd cell_6t
Xbit_r34_c117 bl_117 br_117 wl_34 vdd gnd cell_6t
Xbit_r35_c117 bl_117 br_117 wl_35 vdd gnd cell_6t
Xbit_r36_c117 bl_117 br_117 wl_36 vdd gnd cell_6t
Xbit_r37_c117 bl_117 br_117 wl_37 vdd gnd cell_6t
Xbit_r38_c117 bl_117 br_117 wl_38 vdd gnd cell_6t
Xbit_r39_c117 bl_117 br_117 wl_39 vdd gnd cell_6t
Xbit_r40_c117 bl_117 br_117 wl_40 vdd gnd cell_6t
Xbit_r41_c117 bl_117 br_117 wl_41 vdd gnd cell_6t
Xbit_r42_c117 bl_117 br_117 wl_42 vdd gnd cell_6t
Xbit_r43_c117 bl_117 br_117 wl_43 vdd gnd cell_6t
Xbit_r44_c117 bl_117 br_117 wl_44 vdd gnd cell_6t
Xbit_r45_c117 bl_117 br_117 wl_45 vdd gnd cell_6t
Xbit_r46_c117 bl_117 br_117 wl_46 vdd gnd cell_6t
Xbit_r47_c117 bl_117 br_117 wl_47 vdd gnd cell_6t
Xbit_r48_c117 bl_117 br_117 wl_48 vdd gnd cell_6t
Xbit_r49_c117 bl_117 br_117 wl_49 vdd gnd cell_6t
Xbit_r50_c117 bl_117 br_117 wl_50 vdd gnd cell_6t
Xbit_r51_c117 bl_117 br_117 wl_51 vdd gnd cell_6t
Xbit_r52_c117 bl_117 br_117 wl_52 vdd gnd cell_6t
Xbit_r53_c117 bl_117 br_117 wl_53 vdd gnd cell_6t
Xbit_r54_c117 bl_117 br_117 wl_54 vdd gnd cell_6t
Xbit_r55_c117 bl_117 br_117 wl_55 vdd gnd cell_6t
Xbit_r56_c117 bl_117 br_117 wl_56 vdd gnd cell_6t
Xbit_r57_c117 bl_117 br_117 wl_57 vdd gnd cell_6t
Xbit_r58_c117 bl_117 br_117 wl_58 vdd gnd cell_6t
Xbit_r59_c117 bl_117 br_117 wl_59 vdd gnd cell_6t
Xbit_r60_c117 bl_117 br_117 wl_60 vdd gnd cell_6t
Xbit_r61_c117 bl_117 br_117 wl_61 vdd gnd cell_6t
Xbit_r62_c117 bl_117 br_117 wl_62 vdd gnd cell_6t
Xbit_r63_c117 bl_117 br_117 wl_63 vdd gnd cell_6t
Xbit_r64_c117 bl_117 br_117 wl_64 vdd gnd cell_6t
Xbit_r65_c117 bl_117 br_117 wl_65 vdd gnd cell_6t
Xbit_r66_c117 bl_117 br_117 wl_66 vdd gnd cell_6t
Xbit_r67_c117 bl_117 br_117 wl_67 vdd gnd cell_6t
Xbit_r68_c117 bl_117 br_117 wl_68 vdd gnd cell_6t
Xbit_r69_c117 bl_117 br_117 wl_69 vdd gnd cell_6t
Xbit_r70_c117 bl_117 br_117 wl_70 vdd gnd cell_6t
Xbit_r71_c117 bl_117 br_117 wl_71 vdd gnd cell_6t
Xbit_r72_c117 bl_117 br_117 wl_72 vdd gnd cell_6t
Xbit_r73_c117 bl_117 br_117 wl_73 vdd gnd cell_6t
Xbit_r74_c117 bl_117 br_117 wl_74 vdd gnd cell_6t
Xbit_r75_c117 bl_117 br_117 wl_75 vdd gnd cell_6t
Xbit_r76_c117 bl_117 br_117 wl_76 vdd gnd cell_6t
Xbit_r77_c117 bl_117 br_117 wl_77 vdd gnd cell_6t
Xbit_r78_c117 bl_117 br_117 wl_78 vdd gnd cell_6t
Xbit_r79_c117 bl_117 br_117 wl_79 vdd gnd cell_6t
Xbit_r80_c117 bl_117 br_117 wl_80 vdd gnd cell_6t
Xbit_r81_c117 bl_117 br_117 wl_81 vdd gnd cell_6t
Xbit_r82_c117 bl_117 br_117 wl_82 vdd gnd cell_6t
Xbit_r83_c117 bl_117 br_117 wl_83 vdd gnd cell_6t
Xbit_r84_c117 bl_117 br_117 wl_84 vdd gnd cell_6t
Xbit_r85_c117 bl_117 br_117 wl_85 vdd gnd cell_6t
Xbit_r86_c117 bl_117 br_117 wl_86 vdd gnd cell_6t
Xbit_r87_c117 bl_117 br_117 wl_87 vdd gnd cell_6t
Xbit_r88_c117 bl_117 br_117 wl_88 vdd gnd cell_6t
Xbit_r89_c117 bl_117 br_117 wl_89 vdd gnd cell_6t
Xbit_r90_c117 bl_117 br_117 wl_90 vdd gnd cell_6t
Xbit_r91_c117 bl_117 br_117 wl_91 vdd gnd cell_6t
Xbit_r92_c117 bl_117 br_117 wl_92 vdd gnd cell_6t
Xbit_r93_c117 bl_117 br_117 wl_93 vdd gnd cell_6t
Xbit_r94_c117 bl_117 br_117 wl_94 vdd gnd cell_6t
Xbit_r95_c117 bl_117 br_117 wl_95 vdd gnd cell_6t
Xbit_r96_c117 bl_117 br_117 wl_96 vdd gnd cell_6t
Xbit_r97_c117 bl_117 br_117 wl_97 vdd gnd cell_6t
Xbit_r98_c117 bl_117 br_117 wl_98 vdd gnd cell_6t
Xbit_r99_c117 bl_117 br_117 wl_99 vdd gnd cell_6t
Xbit_r100_c117 bl_117 br_117 wl_100 vdd gnd cell_6t
Xbit_r101_c117 bl_117 br_117 wl_101 vdd gnd cell_6t
Xbit_r102_c117 bl_117 br_117 wl_102 vdd gnd cell_6t
Xbit_r103_c117 bl_117 br_117 wl_103 vdd gnd cell_6t
Xbit_r104_c117 bl_117 br_117 wl_104 vdd gnd cell_6t
Xbit_r105_c117 bl_117 br_117 wl_105 vdd gnd cell_6t
Xbit_r106_c117 bl_117 br_117 wl_106 vdd gnd cell_6t
Xbit_r107_c117 bl_117 br_117 wl_107 vdd gnd cell_6t
Xbit_r108_c117 bl_117 br_117 wl_108 vdd gnd cell_6t
Xbit_r109_c117 bl_117 br_117 wl_109 vdd gnd cell_6t
Xbit_r110_c117 bl_117 br_117 wl_110 vdd gnd cell_6t
Xbit_r111_c117 bl_117 br_117 wl_111 vdd gnd cell_6t
Xbit_r112_c117 bl_117 br_117 wl_112 vdd gnd cell_6t
Xbit_r113_c117 bl_117 br_117 wl_113 vdd gnd cell_6t
Xbit_r114_c117 bl_117 br_117 wl_114 vdd gnd cell_6t
Xbit_r115_c117 bl_117 br_117 wl_115 vdd gnd cell_6t
Xbit_r116_c117 bl_117 br_117 wl_116 vdd gnd cell_6t
Xbit_r117_c117 bl_117 br_117 wl_117 vdd gnd cell_6t
Xbit_r118_c117 bl_117 br_117 wl_118 vdd gnd cell_6t
Xbit_r119_c117 bl_117 br_117 wl_119 vdd gnd cell_6t
Xbit_r120_c117 bl_117 br_117 wl_120 vdd gnd cell_6t
Xbit_r121_c117 bl_117 br_117 wl_121 vdd gnd cell_6t
Xbit_r122_c117 bl_117 br_117 wl_122 vdd gnd cell_6t
Xbit_r123_c117 bl_117 br_117 wl_123 vdd gnd cell_6t
Xbit_r124_c117 bl_117 br_117 wl_124 vdd gnd cell_6t
Xbit_r125_c117 bl_117 br_117 wl_125 vdd gnd cell_6t
Xbit_r126_c117 bl_117 br_117 wl_126 vdd gnd cell_6t
Xbit_r127_c117 bl_117 br_117 wl_127 vdd gnd cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd cell_6t
Xbit_r1_c118 bl_118 br_118 wl_1 vdd gnd cell_6t
Xbit_r2_c118 bl_118 br_118 wl_2 vdd gnd cell_6t
Xbit_r3_c118 bl_118 br_118 wl_3 vdd gnd cell_6t
Xbit_r4_c118 bl_118 br_118 wl_4 vdd gnd cell_6t
Xbit_r5_c118 bl_118 br_118 wl_5 vdd gnd cell_6t
Xbit_r6_c118 bl_118 br_118 wl_6 vdd gnd cell_6t
Xbit_r7_c118 bl_118 br_118 wl_7 vdd gnd cell_6t
Xbit_r8_c118 bl_118 br_118 wl_8 vdd gnd cell_6t
Xbit_r9_c118 bl_118 br_118 wl_9 vdd gnd cell_6t
Xbit_r10_c118 bl_118 br_118 wl_10 vdd gnd cell_6t
Xbit_r11_c118 bl_118 br_118 wl_11 vdd gnd cell_6t
Xbit_r12_c118 bl_118 br_118 wl_12 vdd gnd cell_6t
Xbit_r13_c118 bl_118 br_118 wl_13 vdd gnd cell_6t
Xbit_r14_c118 bl_118 br_118 wl_14 vdd gnd cell_6t
Xbit_r15_c118 bl_118 br_118 wl_15 vdd gnd cell_6t
Xbit_r16_c118 bl_118 br_118 wl_16 vdd gnd cell_6t
Xbit_r17_c118 bl_118 br_118 wl_17 vdd gnd cell_6t
Xbit_r18_c118 bl_118 br_118 wl_18 vdd gnd cell_6t
Xbit_r19_c118 bl_118 br_118 wl_19 vdd gnd cell_6t
Xbit_r20_c118 bl_118 br_118 wl_20 vdd gnd cell_6t
Xbit_r21_c118 bl_118 br_118 wl_21 vdd gnd cell_6t
Xbit_r22_c118 bl_118 br_118 wl_22 vdd gnd cell_6t
Xbit_r23_c118 bl_118 br_118 wl_23 vdd gnd cell_6t
Xbit_r24_c118 bl_118 br_118 wl_24 vdd gnd cell_6t
Xbit_r25_c118 bl_118 br_118 wl_25 vdd gnd cell_6t
Xbit_r26_c118 bl_118 br_118 wl_26 vdd gnd cell_6t
Xbit_r27_c118 bl_118 br_118 wl_27 vdd gnd cell_6t
Xbit_r28_c118 bl_118 br_118 wl_28 vdd gnd cell_6t
Xbit_r29_c118 bl_118 br_118 wl_29 vdd gnd cell_6t
Xbit_r30_c118 bl_118 br_118 wl_30 vdd gnd cell_6t
Xbit_r31_c118 bl_118 br_118 wl_31 vdd gnd cell_6t
Xbit_r32_c118 bl_118 br_118 wl_32 vdd gnd cell_6t
Xbit_r33_c118 bl_118 br_118 wl_33 vdd gnd cell_6t
Xbit_r34_c118 bl_118 br_118 wl_34 vdd gnd cell_6t
Xbit_r35_c118 bl_118 br_118 wl_35 vdd gnd cell_6t
Xbit_r36_c118 bl_118 br_118 wl_36 vdd gnd cell_6t
Xbit_r37_c118 bl_118 br_118 wl_37 vdd gnd cell_6t
Xbit_r38_c118 bl_118 br_118 wl_38 vdd gnd cell_6t
Xbit_r39_c118 bl_118 br_118 wl_39 vdd gnd cell_6t
Xbit_r40_c118 bl_118 br_118 wl_40 vdd gnd cell_6t
Xbit_r41_c118 bl_118 br_118 wl_41 vdd gnd cell_6t
Xbit_r42_c118 bl_118 br_118 wl_42 vdd gnd cell_6t
Xbit_r43_c118 bl_118 br_118 wl_43 vdd gnd cell_6t
Xbit_r44_c118 bl_118 br_118 wl_44 vdd gnd cell_6t
Xbit_r45_c118 bl_118 br_118 wl_45 vdd gnd cell_6t
Xbit_r46_c118 bl_118 br_118 wl_46 vdd gnd cell_6t
Xbit_r47_c118 bl_118 br_118 wl_47 vdd gnd cell_6t
Xbit_r48_c118 bl_118 br_118 wl_48 vdd gnd cell_6t
Xbit_r49_c118 bl_118 br_118 wl_49 vdd gnd cell_6t
Xbit_r50_c118 bl_118 br_118 wl_50 vdd gnd cell_6t
Xbit_r51_c118 bl_118 br_118 wl_51 vdd gnd cell_6t
Xbit_r52_c118 bl_118 br_118 wl_52 vdd gnd cell_6t
Xbit_r53_c118 bl_118 br_118 wl_53 vdd gnd cell_6t
Xbit_r54_c118 bl_118 br_118 wl_54 vdd gnd cell_6t
Xbit_r55_c118 bl_118 br_118 wl_55 vdd gnd cell_6t
Xbit_r56_c118 bl_118 br_118 wl_56 vdd gnd cell_6t
Xbit_r57_c118 bl_118 br_118 wl_57 vdd gnd cell_6t
Xbit_r58_c118 bl_118 br_118 wl_58 vdd gnd cell_6t
Xbit_r59_c118 bl_118 br_118 wl_59 vdd gnd cell_6t
Xbit_r60_c118 bl_118 br_118 wl_60 vdd gnd cell_6t
Xbit_r61_c118 bl_118 br_118 wl_61 vdd gnd cell_6t
Xbit_r62_c118 bl_118 br_118 wl_62 vdd gnd cell_6t
Xbit_r63_c118 bl_118 br_118 wl_63 vdd gnd cell_6t
Xbit_r64_c118 bl_118 br_118 wl_64 vdd gnd cell_6t
Xbit_r65_c118 bl_118 br_118 wl_65 vdd gnd cell_6t
Xbit_r66_c118 bl_118 br_118 wl_66 vdd gnd cell_6t
Xbit_r67_c118 bl_118 br_118 wl_67 vdd gnd cell_6t
Xbit_r68_c118 bl_118 br_118 wl_68 vdd gnd cell_6t
Xbit_r69_c118 bl_118 br_118 wl_69 vdd gnd cell_6t
Xbit_r70_c118 bl_118 br_118 wl_70 vdd gnd cell_6t
Xbit_r71_c118 bl_118 br_118 wl_71 vdd gnd cell_6t
Xbit_r72_c118 bl_118 br_118 wl_72 vdd gnd cell_6t
Xbit_r73_c118 bl_118 br_118 wl_73 vdd gnd cell_6t
Xbit_r74_c118 bl_118 br_118 wl_74 vdd gnd cell_6t
Xbit_r75_c118 bl_118 br_118 wl_75 vdd gnd cell_6t
Xbit_r76_c118 bl_118 br_118 wl_76 vdd gnd cell_6t
Xbit_r77_c118 bl_118 br_118 wl_77 vdd gnd cell_6t
Xbit_r78_c118 bl_118 br_118 wl_78 vdd gnd cell_6t
Xbit_r79_c118 bl_118 br_118 wl_79 vdd gnd cell_6t
Xbit_r80_c118 bl_118 br_118 wl_80 vdd gnd cell_6t
Xbit_r81_c118 bl_118 br_118 wl_81 vdd gnd cell_6t
Xbit_r82_c118 bl_118 br_118 wl_82 vdd gnd cell_6t
Xbit_r83_c118 bl_118 br_118 wl_83 vdd gnd cell_6t
Xbit_r84_c118 bl_118 br_118 wl_84 vdd gnd cell_6t
Xbit_r85_c118 bl_118 br_118 wl_85 vdd gnd cell_6t
Xbit_r86_c118 bl_118 br_118 wl_86 vdd gnd cell_6t
Xbit_r87_c118 bl_118 br_118 wl_87 vdd gnd cell_6t
Xbit_r88_c118 bl_118 br_118 wl_88 vdd gnd cell_6t
Xbit_r89_c118 bl_118 br_118 wl_89 vdd gnd cell_6t
Xbit_r90_c118 bl_118 br_118 wl_90 vdd gnd cell_6t
Xbit_r91_c118 bl_118 br_118 wl_91 vdd gnd cell_6t
Xbit_r92_c118 bl_118 br_118 wl_92 vdd gnd cell_6t
Xbit_r93_c118 bl_118 br_118 wl_93 vdd gnd cell_6t
Xbit_r94_c118 bl_118 br_118 wl_94 vdd gnd cell_6t
Xbit_r95_c118 bl_118 br_118 wl_95 vdd gnd cell_6t
Xbit_r96_c118 bl_118 br_118 wl_96 vdd gnd cell_6t
Xbit_r97_c118 bl_118 br_118 wl_97 vdd gnd cell_6t
Xbit_r98_c118 bl_118 br_118 wl_98 vdd gnd cell_6t
Xbit_r99_c118 bl_118 br_118 wl_99 vdd gnd cell_6t
Xbit_r100_c118 bl_118 br_118 wl_100 vdd gnd cell_6t
Xbit_r101_c118 bl_118 br_118 wl_101 vdd gnd cell_6t
Xbit_r102_c118 bl_118 br_118 wl_102 vdd gnd cell_6t
Xbit_r103_c118 bl_118 br_118 wl_103 vdd gnd cell_6t
Xbit_r104_c118 bl_118 br_118 wl_104 vdd gnd cell_6t
Xbit_r105_c118 bl_118 br_118 wl_105 vdd gnd cell_6t
Xbit_r106_c118 bl_118 br_118 wl_106 vdd gnd cell_6t
Xbit_r107_c118 bl_118 br_118 wl_107 vdd gnd cell_6t
Xbit_r108_c118 bl_118 br_118 wl_108 vdd gnd cell_6t
Xbit_r109_c118 bl_118 br_118 wl_109 vdd gnd cell_6t
Xbit_r110_c118 bl_118 br_118 wl_110 vdd gnd cell_6t
Xbit_r111_c118 bl_118 br_118 wl_111 vdd gnd cell_6t
Xbit_r112_c118 bl_118 br_118 wl_112 vdd gnd cell_6t
Xbit_r113_c118 bl_118 br_118 wl_113 vdd gnd cell_6t
Xbit_r114_c118 bl_118 br_118 wl_114 vdd gnd cell_6t
Xbit_r115_c118 bl_118 br_118 wl_115 vdd gnd cell_6t
Xbit_r116_c118 bl_118 br_118 wl_116 vdd gnd cell_6t
Xbit_r117_c118 bl_118 br_118 wl_117 vdd gnd cell_6t
Xbit_r118_c118 bl_118 br_118 wl_118 vdd gnd cell_6t
Xbit_r119_c118 bl_118 br_118 wl_119 vdd gnd cell_6t
Xbit_r120_c118 bl_118 br_118 wl_120 vdd gnd cell_6t
Xbit_r121_c118 bl_118 br_118 wl_121 vdd gnd cell_6t
Xbit_r122_c118 bl_118 br_118 wl_122 vdd gnd cell_6t
Xbit_r123_c118 bl_118 br_118 wl_123 vdd gnd cell_6t
Xbit_r124_c118 bl_118 br_118 wl_124 vdd gnd cell_6t
Xbit_r125_c118 bl_118 br_118 wl_125 vdd gnd cell_6t
Xbit_r126_c118 bl_118 br_118 wl_126 vdd gnd cell_6t
Xbit_r127_c118 bl_118 br_118 wl_127 vdd gnd cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd cell_6t
Xbit_r1_c119 bl_119 br_119 wl_1 vdd gnd cell_6t
Xbit_r2_c119 bl_119 br_119 wl_2 vdd gnd cell_6t
Xbit_r3_c119 bl_119 br_119 wl_3 vdd gnd cell_6t
Xbit_r4_c119 bl_119 br_119 wl_4 vdd gnd cell_6t
Xbit_r5_c119 bl_119 br_119 wl_5 vdd gnd cell_6t
Xbit_r6_c119 bl_119 br_119 wl_6 vdd gnd cell_6t
Xbit_r7_c119 bl_119 br_119 wl_7 vdd gnd cell_6t
Xbit_r8_c119 bl_119 br_119 wl_8 vdd gnd cell_6t
Xbit_r9_c119 bl_119 br_119 wl_9 vdd gnd cell_6t
Xbit_r10_c119 bl_119 br_119 wl_10 vdd gnd cell_6t
Xbit_r11_c119 bl_119 br_119 wl_11 vdd gnd cell_6t
Xbit_r12_c119 bl_119 br_119 wl_12 vdd gnd cell_6t
Xbit_r13_c119 bl_119 br_119 wl_13 vdd gnd cell_6t
Xbit_r14_c119 bl_119 br_119 wl_14 vdd gnd cell_6t
Xbit_r15_c119 bl_119 br_119 wl_15 vdd gnd cell_6t
Xbit_r16_c119 bl_119 br_119 wl_16 vdd gnd cell_6t
Xbit_r17_c119 bl_119 br_119 wl_17 vdd gnd cell_6t
Xbit_r18_c119 bl_119 br_119 wl_18 vdd gnd cell_6t
Xbit_r19_c119 bl_119 br_119 wl_19 vdd gnd cell_6t
Xbit_r20_c119 bl_119 br_119 wl_20 vdd gnd cell_6t
Xbit_r21_c119 bl_119 br_119 wl_21 vdd gnd cell_6t
Xbit_r22_c119 bl_119 br_119 wl_22 vdd gnd cell_6t
Xbit_r23_c119 bl_119 br_119 wl_23 vdd gnd cell_6t
Xbit_r24_c119 bl_119 br_119 wl_24 vdd gnd cell_6t
Xbit_r25_c119 bl_119 br_119 wl_25 vdd gnd cell_6t
Xbit_r26_c119 bl_119 br_119 wl_26 vdd gnd cell_6t
Xbit_r27_c119 bl_119 br_119 wl_27 vdd gnd cell_6t
Xbit_r28_c119 bl_119 br_119 wl_28 vdd gnd cell_6t
Xbit_r29_c119 bl_119 br_119 wl_29 vdd gnd cell_6t
Xbit_r30_c119 bl_119 br_119 wl_30 vdd gnd cell_6t
Xbit_r31_c119 bl_119 br_119 wl_31 vdd gnd cell_6t
Xbit_r32_c119 bl_119 br_119 wl_32 vdd gnd cell_6t
Xbit_r33_c119 bl_119 br_119 wl_33 vdd gnd cell_6t
Xbit_r34_c119 bl_119 br_119 wl_34 vdd gnd cell_6t
Xbit_r35_c119 bl_119 br_119 wl_35 vdd gnd cell_6t
Xbit_r36_c119 bl_119 br_119 wl_36 vdd gnd cell_6t
Xbit_r37_c119 bl_119 br_119 wl_37 vdd gnd cell_6t
Xbit_r38_c119 bl_119 br_119 wl_38 vdd gnd cell_6t
Xbit_r39_c119 bl_119 br_119 wl_39 vdd gnd cell_6t
Xbit_r40_c119 bl_119 br_119 wl_40 vdd gnd cell_6t
Xbit_r41_c119 bl_119 br_119 wl_41 vdd gnd cell_6t
Xbit_r42_c119 bl_119 br_119 wl_42 vdd gnd cell_6t
Xbit_r43_c119 bl_119 br_119 wl_43 vdd gnd cell_6t
Xbit_r44_c119 bl_119 br_119 wl_44 vdd gnd cell_6t
Xbit_r45_c119 bl_119 br_119 wl_45 vdd gnd cell_6t
Xbit_r46_c119 bl_119 br_119 wl_46 vdd gnd cell_6t
Xbit_r47_c119 bl_119 br_119 wl_47 vdd gnd cell_6t
Xbit_r48_c119 bl_119 br_119 wl_48 vdd gnd cell_6t
Xbit_r49_c119 bl_119 br_119 wl_49 vdd gnd cell_6t
Xbit_r50_c119 bl_119 br_119 wl_50 vdd gnd cell_6t
Xbit_r51_c119 bl_119 br_119 wl_51 vdd gnd cell_6t
Xbit_r52_c119 bl_119 br_119 wl_52 vdd gnd cell_6t
Xbit_r53_c119 bl_119 br_119 wl_53 vdd gnd cell_6t
Xbit_r54_c119 bl_119 br_119 wl_54 vdd gnd cell_6t
Xbit_r55_c119 bl_119 br_119 wl_55 vdd gnd cell_6t
Xbit_r56_c119 bl_119 br_119 wl_56 vdd gnd cell_6t
Xbit_r57_c119 bl_119 br_119 wl_57 vdd gnd cell_6t
Xbit_r58_c119 bl_119 br_119 wl_58 vdd gnd cell_6t
Xbit_r59_c119 bl_119 br_119 wl_59 vdd gnd cell_6t
Xbit_r60_c119 bl_119 br_119 wl_60 vdd gnd cell_6t
Xbit_r61_c119 bl_119 br_119 wl_61 vdd gnd cell_6t
Xbit_r62_c119 bl_119 br_119 wl_62 vdd gnd cell_6t
Xbit_r63_c119 bl_119 br_119 wl_63 vdd gnd cell_6t
Xbit_r64_c119 bl_119 br_119 wl_64 vdd gnd cell_6t
Xbit_r65_c119 bl_119 br_119 wl_65 vdd gnd cell_6t
Xbit_r66_c119 bl_119 br_119 wl_66 vdd gnd cell_6t
Xbit_r67_c119 bl_119 br_119 wl_67 vdd gnd cell_6t
Xbit_r68_c119 bl_119 br_119 wl_68 vdd gnd cell_6t
Xbit_r69_c119 bl_119 br_119 wl_69 vdd gnd cell_6t
Xbit_r70_c119 bl_119 br_119 wl_70 vdd gnd cell_6t
Xbit_r71_c119 bl_119 br_119 wl_71 vdd gnd cell_6t
Xbit_r72_c119 bl_119 br_119 wl_72 vdd gnd cell_6t
Xbit_r73_c119 bl_119 br_119 wl_73 vdd gnd cell_6t
Xbit_r74_c119 bl_119 br_119 wl_74 vdd gnd cell_6t
Xbit_r75_c119 bl_119 br_119 wl_75 vdd gnd cell_6t
Xbit_r76_c119 bl_119 br_119 wl_76 vdd gnd cell_6t
Xbit_r77_c119 bl_119 br_119 wl_77 vdd gnd cell_6t
Xbit_r78_c119 bl_119 br_119 wl_78 vdd gnd cell_6t
Xbit_r79_c119 bl_119 br_119 wl_79 vdd gnd cell_6t
Xbit_r80_c119 bl_119 br_119 wl_80 vdd gnd cell_6t
Xbit_r81_c119 bl_119 br_119 wl_81 vdd gnd cell_6t
Xbit_r82_c119 bl_119 br_119 wl_82 vdd gnd cell_6t
Xbit_r83_c119 bl_119 br_119 wl_83 vdd gnd cell_6t
Xbit_r84_c119 bl_119 br_119 wl_84 vdd gnd cell_6t
Xbit_r85_c119 bl_119 br_119 wl_85 vdd gnd cell_6t
Xbit_r86_c119 bl_119 br_119 wl_86 vdd gnd cell_6t
Xbit_r87_c119 bl_119 br_119 wl_87 vdd gnd cell_6t
Xbit_r88_c119 bl_119 br_119 wl_88 vdd gnd cell_6t
Xbit_r89_c119 bl_119 br_119 wl_89 vdd gnd cell_6t
Xbit_r90_c119 bl_119 br_119 wl_90 vdd gnd cell_6t
Xbit_r91_c119 bl_119 br_119 wl_91 vdd gnd cell_6t
Xbit_r92_c119 bl_119 br_119 wl_92 vdd gnd cell_6t
Xbit_r93_c119 bl_119 br_119 wl_93 vdd gnd cell_6t
Xbit_r94_c119 bl_119 br_119 wl_94 vdd gnd cell_6t
Xbit_r95_c119 bl_119 br_119 wl_95 vdd gnd cell_6t
Xbit_r96_c119 bl_119 br_119 wl_96 vdd gnd cell_6t
Xbit_r97_c119 bl_119 br_119 wl_97 vdd gnd cell_6t
Xbit_r98_c119 bl_119 br_119 wl_98 vdd gnd cell_6t
Xbit_r99_c119 bl_119 br_119 wl_99 vdd gnd cell_6t
Xbit_r100_c119 bl_119 br_119 wl_100 vdd gnd cell_6t
Xbit_r101_c119 bl_119 br_119 wl_101 vdd gnd cell_6t
Xbit_r102_c119 bl_119 br_119 wl_102 vdd gnd cell_6t
Xbit_r103_c119 bl_119 br_119 wl_103 vdd gnd cell_6t
Xbit_r104_c119 bl_119 br_119 wl_104 vdd gnd cell_6t
Xbit_r105_c119 bl_119 br_119 wl_105 vdd gnd cell_6t
Xbit_r106_c119 bl_119 br_119 wl_106 vdd gnd cell_6t
Xbit_r107_c119 bl_119 br_119 wl_107 vdd gnd cell_6t
Xbit_r108_c119 bl_119 br_119 wl_108 vdd gnd cell_6t
Xbit_r109_c119 bl_119 br_119 wl_109 vdd gnd cell_6t
Xbit_r110_c119 bl_119 br_119 wl_110 vdd gnd cell_6t
Xbit_r111_c119 bl_119 br_119 wl_111 vdd gnd cell_6t
Xbit_r112_c119 bl_119 br_119 wl_112 vdd gnd cell_6t
Xbit_r113_c119 bl_119 br_119 wl_113 vdd gnd cell_6t
Xbit_r114_c119 bl_119 br_119 wl_114 vdd gnd cell_6t
Xbit_r115_c119 bl_119 br_119 wl_115 vdd gnd cell_6t
Xbit_r116_c119 bl_119 br_119 wl_116 vdd gnd cell_6t
Xbit_r117_c119 bl_119 br_119 wl_117 vdd gnd cell_6t
Xbit_r118_c119 bl_119 br_119 wl_118 vdd gnd cell_6t
Xbit_r119_c119 bl_119 br_119 wl_119 vdd gnd cell_6t
Xbit_r120_c119 bl_119 br_119 wl_120 vdd gnd cell_6t
Xbit_r121_c119 bl_119 br_119 wl_121 vdd gnd cell_6t
Xbit_r122_c119 bl_119 br_119 wl_122 vdd gnd cell_6t
Xbit_r123_c119 bl_119 br_119 wl_123 vdd gnd cell_6t
Xbit_r124_c119 bl_119 br_119 wl_124 vdd gnd cell_6t
Xbit_r125_c119 bl_119 br_119 wl_125 vdd gnd cell_6t
Xbit_r126_c119 bl_119 br_119 wl_126 vdd gnd cell_6t
Xbit_r127_c119 bl_119 br_119 wl_127 vdd gnd cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd cell_6t
Xbit_r1_c120 bl_120 br_120 wl_1 vdd gnd cell_6t
Xbit_r2_c120 bl_120 br_120 wl_2 vdd gnd cell_6t
Xbit_r3_c120 bl_120 br_120 wl_3 vdd gnd cell_6t
Xbit_r4_c120 bl_120 br_120 wl_4 vdd gnd cell_6t
Xbit_r5_c120 bl_120 br_120 wl_5 vdd gnd cell_6t
Xbit_r6_c120 bl_120 br_120 wl_6 vdd gnd cell_6t
Xbit_r7_c120 bl_120 br_120 wl_7 vdd gnd cell_6t
Xbit_r8_c120 bl_120 br_120 wl_8 vdd gnd cell_6t
Xbit_r9_c120 bl_120 br_120 wl_9 vdd gnd cell_6t
Xbit_r10_c120 bl_120 br_120 wl_10 vdd gnd cell_6t
Xbit_r11_c120 bl_120 br_120 wl_11 vdd gnd cell_6t
Xbit_r12_c120 bl_120 br_120 wl_12 vdd gnd cell_6t
Xbit_r13_c120 bl_120 br_120 wl_13 vdd gnd cell_6t
Xbit_r14_c120 bl_120 br_120 wl_14 vdd gnd cell_6t
Xbit_r15_c120 bl_120 br_120 wl_15 vdd gnd cell_6t
Xbit_r16_c120 bl_120 br_120 wl_16 vdd gnd cell_6t
Xbit_r17_c120 bl_120 br_120 wl_17 vdd gnd cell_6t
Xbit_r18_c120 bl_120 br_120 wl_18 vdd gnd cell_6t
Xbit_r19_c120 bl_120 br_120 wl_19 vdd gnd cell_6t
Xbit_r20_c120 bl_120 br_120 wl_20 vdd gnd cell_6t
Xbit_r21_c120 bl_120 br_120 wl_21 vdd gnd cell_6t
Xbit_r22_c120 bl_120 br_120 wl_22 vdd gnd cell_6t
Xbit_r23_c120 bl_120 br_120 wl_23 vdd gnd cell_6t
Xbit_r24_c120 bl_120 br_120 wl_24 vdd gnd cell_6t
Xbit_r25_c120 bl_120 br_120 wl_25 vdd gnd cell_6t
Xbit_r26_c120 bl_120 br_120 wl_26 vdd gnd cell_6t
Xbit_r27_c120 bl_120 br_120 wl_27 vdd gnd cell_6t
Xbit_r28_c120 bl_120 br_120 wl_28 vdd gnd cell_6t
Xbit_r29_c120 bl_120 br_120 wl_29 vdd gnd cell_6t
Xbit_r30_c120 bl_120 br_120 wl_30 vdd gnd cell_6t
Xbit_r31_c120 bl_120 br_120 wl_31 vdd gnd cell_6t
Xbit_r32_c120 bl_120 br_120 wl_32 vdd gnd cell_6t
Xbit_r33_c120 bl_120 br_120 wl_33 vdd gnd cell_6t
Xbit_r34_c120 bl_120 br_120 wl_34 vdd gnd cell_6t
Xbit_r35_c120 bl_120 br_120 wl_35 vdd gnd cell_6t
Xbit_r36_c120 bl_120 br_120 wl_36 vdd gnd cell_6t
Xbit_r37_c120 bl_120 br_120 wl_37 vdd gnd cell_6t
Xbit_r38_c120 bl_120 br_120 wl_38 vdd gnd cell_6t
Xbit_r39_c120 bl_120 br_120 wl_39 vdd gnd cell_6t
Xbit_r40_c120 bl_120 br_120 wl_40 vdd gnd cell_6t
Xbit_r41_c120 bl_120 br_120 wl_41 vdd gnd cell_6t
Xbit_r42_c120 bl_120 br_120 wl_42 vdd gnd cell_6t
Xbit_r43_c120 bl_120 br_120 wl_43 vdd gnd cell_6t
Xbit_r44_c120 bl_120 br_120 wl_44 vdd gnd cell_6t
Xbit_r45_c120 bl_120 br_120 wl_45 vdd gnd cell_6t
Xbit_r46_c120 bl_120 br_120 wl_46 vdd gnd cell_6t
Xbit_r47_c120 bl_120 br_120 wl_47 vdd gnd cell_6t
Xbit_r48_c120 bl_120 br_120 wl_48 vdd gnd cell_6t
Xbit_r49_c120 bl_120 br_120 wl_49 vdd gnd cell_6t
Xbit_r50_c120 bl_120 br_120 wl_50 vdd gnd cell_6t
Xbit_r51_c120 bl_120 br_120 wl_51 vdd gnd cell_6t
Xbit_r52_c120 bl_120 br_120 wl_52 vdd gnd cell_6t
Xbit_r53_c120 bl_120 br_120 wl_53 vdd gnd cell_6t
Xbit_r54_c120 bl_120 br_120 wl_54 vdd gnd cell_6t
Xbit_r55_c120 bl_120 br_120 wl_55 vdd gnd cell_6t
Xbit_r56_c120 bl_120 br_120 wl_56 vdd gnd cell_6t
Xbit_r57_c120 bl_120 br_120 wl_57 vdd gnd cell_6t
Xbit_r58_c120 bl_120 br_120 wl_58 vdd gnd cell_6t
Xbit_r59_c120 bl_120 br_120 wl_59 vdd gnd cell_6t
Xbit_r60_c120 bl_120 br_120 wl_60 vdd gnd cell_6t
Xbit_r61_c120 bl_120 br_120 wl_61 vdd gnd cell_6t
Xbit_r62_c120 bl_120 br_120 wl_62 vdd gnd cell_6t
Xbit_r63_c120 bl_120 br_120 wl_63 vdd gnd cell_6t
Xbit_r64_c120 bl_120 br_120 wl_64 vdd gnd cell_6t
Xbit_r65_c120 bl_120 br_120 wl_65 vdd gnd cell_6t
Xbit_r66_c120 bl_120 br_120 wl_66 vdd gnd cell_6t
Xbit_r67_c120 bl_120 br_120 wl_67 vdd gnd cell_6t
Xbit_r68_c120 bl_120 br_120 wl_68 vdd gnd cell_6t
Xbit_r69_c120 bl_120 br_120 wl_69 vdd gnd cell_6t
Xbit_r70_c120 bl_120 br_120 wl_70 vdd gnd cell_6t
Xbit_r71_c120 bl_120 br_120 wl_71 vdd gnd cell_6t
Xbit_r72_c120 bl_120 br_120 wl_72 vdd gnd cell_6t
Xbit_r73_c120 bl_120 br_120 wl_73 vdd gnd cell_6t
Xbit_r74_c120 bl_120 br_120 wl_74 vdd gnd cell_6t
Xbit_r75_c120 bl_120 br_120 wl_75 vdd gnd cell_6t
Xbit_r76_c120 bl_120 br_120 wl_76 vdd gnd cell_6t
Xbit_r77_c120 bl_120 br_120 wl_77 vdd gnd cell_6t
Xbit_r78_c120 bl_120 br_120 wl_78 vdd gnd cell_6t
Xbit_r79_c120 bl_120 br_120 wl_79 vdd gnd cell_6t
Xbit_r80_c120 bl_120 br_120 wl_80 vdd gnd cell_6t
Xbit_r81_c120 bl_120 br_120 wl_81 vdd gnd cell_6t
Xbit_r82_c120 bl_120 br_120 wl_82 vdd gnd cell_6t
Xbit_r83_c120 bl_120 br_120 wl_83 vdd gnd cell_6t
Xbit_r84_c120 bl_120 br_120 wl_84 vdd gnd cell_6t
Xbit_r85_c120 bl_120 br_120 wl_85 vdd gnd cell_6t
Xbit_r86_c120 bl_120 br_120 wl_86 vdd gnd cell_6t
Xbit_r87_c120 bl_120 br_120 wl_87 vdd gnd cell_6t
Xbit_r88_c120 bl_120 br_120 wl_88 vdd gnd cell_6t
Xbit_r89_c120 bl_120 br_120 wl_89 vdd gnd cell_6t
Xbit_r90_c120 bl_120 br_120 wl_90 vdd gnd cell_6t
Xbit_r91_c120 bl_120 br_120 wl_91 vdd gnd cell_6t
Xbit_r92_c120 bl_120 br_120 wl_92 vdd gnd cell_6t
Xbit_r93_c120 bl_120 br_120 wl_93 vdd gnd cell_6t
Xbit_r94_c120 bl_120 br_120 wl_94 vdd gnd cell_6t
Xbit_r95_c120 bl_120 br_120 wl_95 vdd gnd cell_6t
Xbit_r96_c120 bl_120 br_120 wl_96 vdd gnd cell_6t
Xbit_r97_c120 bl_120 br_120 wl_97 vdd gnd cell_6t
Xbit_r98_c120 bl_120 br_120 wl_98 vdd gnd cell_6t
Xbit_r99_c120 bl_120 br_120 wl_99 vdd gnd cell_6t
Xbit_r100_c120 bl_120 br_120 wl_100 vdd gnd cell_6t
Xbit_r101_c120 bl_120 br_120 wl_101 vdd gnd cell_6t
Xbit_r102_c120 bl_120 br_120 wl_102 vdd gnd cell_6t
Xbit_r103_c120 bl_120 br_120 wl_103 vdd gnd cell_6t
Xbit_r104_c120 bl_120 br_120 wl_104 vdd gnd cell_6t
Xbit_r105_c120 bl_120 br_120 wl_105 vdd gnd cell_6t
Xbit_r106_c120 bl_120 br_120 wl_106 vdd gnd cell_6t
Xbit_r107_c120 bl_120 br_120 wl_107 vdd gnd cell_6t
Xbit_r108_c120 bl_120 br_120 wl_108 vdd gnd cell_6t
Xbit_r109_c120 bl_120 br_120 wl_109 vdd gnd cell_6t
Xbit_r110_c120 bl_120 br_120 wl_110 vdd gnd cell_6t
Xbit_r111_c120 bl_120 br_120 wl_111 vdd gnd cell_6t
Xbit_r112_c120 bl_120 br_120 wl_112 vdd gnd cell_6t
Xbit_r113_c120 bl_120 br_120 wl_113 vdd gnd cell_6t
Xbit_r114_c120 bl_120 br_120 wl_114 vdd gnd cell_6t
Xbit_r115_c120 bl_120 br_120 wl_115 vdd gnd cell_6t
Xbit_r116_c120 bl_120 br_120 wl_116 vdd gnd cell_6t
Xbit_r117_c120 bl_120 br_120 wl_117 vdd gnd cell_6t
Xbit_r118_c120 bl_120 br_120 wl_118 vdd gnd cell_6t
Xbit_r119_c120 bl_120 br_120 wl_119 vdd gnd cell_6t
Xbit_r120_c120 bl_120 br_120 wl_120 vdd gnd cell_6t
Xbit_r121_c120 bl_120 br_120 wl_121 vdd gnd cell_6t
Xbit_r122_c120 bl_120 br_120 wl_122 vdd gnd cell_6t
Xbit_r123_c120 bl_120 br_120 wl_123 vdd gnd cell_6t
Xbit_r124_c120 bl_120 br_120 wl_124 vdd gnd cell_6t
Xbit_r125_c120 bl_120 br_120 wl_125 vdd gnd cell_6t
Xbit_r126_c120 bl_120 br_120 wl_126 vdd gnd cell_6t
Xbit_r127_c120 bl_120 br_120 wl_127 vdd gnd cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd cell_6t
Xbit_r1_c121 bl_121 br_121 wl_1 vdd gnd cell_6t
Xbit_r2_c121 bl_121 br_121 wl_2 vdd gnd cell_6t
Xbit_r3_c121 bl_121 br_121 wl_3 vdd gnd cell_6t
Xbit_r4_c121 bl_121 br_121 wl_4 vdd gnd cell_6t
Xbit_r5_c121 bl_121 br_121 wl_5 vdd gnd cell_6t
Xbit_r6_c121 bl_121 br_121 wl_6 vdd gnd cell_6t
Xbit_r7_c121 bl_121 br_121 wl_7 vdd gnd cell_6t
Xbit_r8_c121 bl_121 br_121 wl_8 vdd gnd cell_6t
Xbit_r9_c121 bl_121 br_121 wl_9 vdd gnd cell_6t
Xbit_r10_c121 bl_121 br_121 wl_10 vdd gnd cell_6t
Xbit_r11_c121 bl_121 br_121 wl_11 vdd gnd cell_6t
Xbit_r12_c121 bl_121 br_121 wl_12 vdd gnd cell_6t
Xbit_r13_c121 bl_121 br_121 wl_13 vdd gnd cell_6t
Xbit_r14_c121 bl_121 br_121 wl_14 vdd gnd cell_6t
Xbit_r15_c121 bl_121 br_121 wl_15 vdd gnd cell_6t
Xbit_r16_c121 bl_121 br_121 wl_16 vdd gnd cell_6t
Xbit_r17_c121 bl_121 br_121 wl_17 vdd gnd cell_6t
Xbit_r18_c121 bl_121 br_121 wl_18 vdd gnd cell_6t
Xbit_r19_c121 bl_121 br_121 wl_19 vdd gnd cell_6t
Xbit_r20_c121 bl_121 br_121 wl_20 vdd gnd cell_6t
Xbit_r21_c121 bl_121 br_121 wl_21 vdd gnd cell_6t
Xbit_r22_c121 bl_121 br_121 wl_22 vdd gnd cell_6t
Xbit_r23_c121 bl_121 br_121 wl_23 vdd gnd cell_6t
Xbit_r24_c121 bl_121 br_121 wl_24 vdd gnd cell_6t
Xbit_r25_c121 bl_121 br_121 wl_25 vdd gnd cell_6t
Xbit_r26_c121 bl_121 br_121 wl_26 vdd gnd cell_6t
Xbit_r27_c121 bl_121 br_121 wl_27 vdd gnd cell_6t
Xbit_r28_c121 bl_121 br_121 wl_28 vdd gnd cell_6t
Xbit_r29_c121 bl_121 br_121 wl_29 vdd gnd cell_6t
Xbit_r30_c121 bl_121 br_121 wl_30 vdd gnd cell_6t
Xbit_r31_c121 bl_121 br_121 wl_31 vdd gnd cell_6t
Xbit_r32_c121 bl_121 br_121 wl_32 vdd gnd cell_6t
Xbit_r33_c121 bl_121 br_121 wl_33 vdd gnd cell_6t
Xbit_r34_c121 bl_121 br_121 wl_34 vdd gnd cell_6t
Xbit_r35_c121 bl_121 br_121 wl_35 vdd gnd cell_6t
Xbit_r36_c121 bl_121 br_121 wl_36 vdd gnd cell_6t
Xbit_r37_c121 bl_121 br_121 wl_37 vdd gnd cell_6t
Xbit_r38_c121 bl_121 br_121 wl_38 vdd gnd cell_6t
Xbit_r39_c121 bl_121 br_121 wl_39 vdd gnd cell_6t
Xbit_r40_c121 bl_121 br_121 wl_40 vdd gnd cell_6t
Xbit_r41_c121 bl_121 br_121 wl_41 vdd gnd cell_6t
Xbit_r42_c121 bl_121 br_121 wl_42 vdd gnd cell_6t
Xbit_r43_c121 bl_121 br_121 wl_43 vdd gnd cell_6t
Xbit_r44_c121 bl_121 br_121 wl_44 vdd gnd cell_6t
Xbit_r45_c121 bl_121 br_121 wl_45 vdd gnd cell_6t
Xbit_r46_c121 bl_121 br_121 wl_46 vdd gnd cell_6t
Xbit_r47_c121 bl_121 br_121 wl_47 vdd gnd cell_6t
Xbit_r48_c121 bl_121 br_121 wl_48 vdd gnd cell_6t
Xbit_r49_c121 bl_121 br_121 wl_49 vdd gnd cell_6t
Xbit_r50_c121 bl_121 br_121 wl_50 vdd gnd cell_6t
Xbit_r51_c121 bl_121 br_121 wl_51 vdd gnd cell_6t
Xbit_r52_c121 bl_121 br_121 wl_52 vdd gnd cell_6t
Xbit_r53_c121 bl_121 br_121 wl_53 vdd gnd cell_6t
Xbit_r54_c121 bl_121 br_121 wl_54 vdd gnd cell_6t
Xbit_r55_c121 bl_121 br_121 wl_55 vdd gnd cell_6t
Xbit_r56_c121 bl_121 br_121 wl_56 vdd gnd cell_6t
Xbit_r57_c121 bl_121 br_121 wl_57 vdd gnd cell_6t
Xbit_r58_c121 bl_121 br_121 wl_58 vdd gnd cell_6t
Xbit_r59_c121 bl_121 br_121 wl_59 vdd gnd cell_6t
Xbit_r60_c121 bl_121 br_121 wl_60 vdd gnd cell_6t
Xbit_r61_c121 bl_121 br_121 wl_61 vdd gnd cell_6t
Xbit_r62_c121 bl_121 br_121 wl_62 vdd gnd cell_6t
Xbit_r63_c121 bl_121 br_121 wl_63 vdd gnd cell_6t
Xbit_r64_c121 bl_121 br_121 wl_64 vdd gnd cell_6t
Xbit_r65_c121 bl_121 br_121 wl_65 vdd gnd cell_6t
Xbit_r66_c121 bl_121 br_121 wl_66 vdd gnd cell_6t
Xbit_r67_c121 bl_121 br_121 wl_67 vdd gnd cell_6t
Xbit_r68_c121 bl_121 br_121 wl_68 vdd gnd cell_6t
Xbit_r69_c121 bl_121 br_121 wl_69 vdd gnd cell_6t
Xbit_r70_c121 bl_121 br_121 wl_70 vdd gnd cell_6t
Xbit_r71_c121 bl_121 br_121 wl_71 vdd gnd cell_6t
Xbit_r72_c121 bl_121 br_121 wl_72 vdd gnd cell_6t
Xbit_r73_c121 bl_121 br_121 wl_73 vdd gnd cell_6t
Xbit_r74_c121 bl_121 br_121 wl_74 vdd gnd cell_6t
Xbit_r75_c121 bl_121 br_121 wl_75 vdd gnd cell_6t
Xbit_r76_c121 bl_121 br_121 wl_76 vdd gnd cell_6t
Xbit_r77_c121 bl_121 br_121 wl_77 vdd gnd cell_6t
Xbit_r78_c121 bl_121 br_121 wl_78 vdd gnd cell_6t
Xbit_r79_c121 bl_121 br_121 wl_79 vdd gnd cell_6t
Xbit_r80_c121 bl_121 br_121 wl_80 vdd gnd cell_6t
Xbit_r81_c121 bl_121 br_121 wl_81 vdd gnd cell_6t
Xbit_r82_c121 bl_121 br_121 wl_82 vdd gnd cell_6t
Xbit_r83_c121 bl_121 br_121 wl_83 vdd gnd cell_6t
Xbit_r84_c121 bl_121 br_121 wl_84 vdd gnd cell_6t
Xbit_r85_c121 bl_121 br_121 wl_85 vdd gnd cell_6t
Xbit_r86_c121 bl_121 br_121 wl_86 vdd gnd cell_6t
Xbit_r87_c121 bl_121 br_121 wl_87 vdd gnd cell_6t
Xbit_r88_c121 bl_121 br_121 wl_88 vdd gnd cell_6t
Xbit_r89_c121 bl_121 br_121 wl_89 vdd gnd cell_6t
Xbit_r90_c121 bl_121 br_121 wl_90 vdd gnd cell_6t
Xbit_r91_c121 bl_121 br_121 wl_91 vdd gnd cell_6t
Xbit_r92_c121 bl_121 br_121 wl_92 vdd gnd cell_6t
Xbit_r93_c121 bl_121 br_121 wl_93 vdd gnd cell_6t
Xbit_r94_c121 bl_121 br_121 wl_94 vdd gnd cell_6t
Xbit_r95_c121 bl_121 br_121 wl_95 vdd gnd cell_6t
Xbit_r96_c121 bl_121 br_121 wl_96 vdd gnd cell_6t
Xbit_r97_c121 bl_121 br_121 wl_97 vdd gnd cell_6t
Xbit_r98_c121 bl_121 br_121 wl_98 vdd gnd cell_6t
Xbit_r99_c121 bl_121 br_121 wl_99 vdd gnd cell_6t
Xbit_r100_c121 bl_121 br_121 wl_100 vdd gnd cell_6t
Xbit_r101_c121 bl_121 br_121 wl_101 vdd gnd cell_6t
Xbit_r102_c121 bl_121 br_121 wl_102 vdd gnd cell_6t
Xbit_r103_c121 bl_121 br_121 wl_103 vdd gnd cell_6t
Xbit_r104_c121 bl_121 br_121 wl_104 vdd gnd cell_6t
Xbit_r105_c121 bl_121 br_121 wl_105 vdd gnd cell_6t
Xbit_r106_c121 bl_121 br_121 wl_106 vdd gnd cell_6t
Xbit_r107_c121 bl_121 br_121 wl_107 vdd gnd cell_6t
Xbit_r108_c121 bl_121 br_121 wl_108 vdd gnd cell_6t
Xbit_r109_c121 bl_121 br_121 wl_109 vdd gnd cell_6t
Xbit_r110_c121 bl_121 br_121 wl_110 vdd gnd cell_6t
Xbit_r111_c121 bl_121 br_121 wl_111 vdd gnd cell_6t
Xbit_r112_c121 bl_121 br_121 wl_112 vdd gnd cell_6t
Xbit_r113_c121 bl_121 br_121 wl_113 vdd gnd cell_6t
Xbit_r114_c121 bl_121 br_121 wl_114 vdd gnd cell_6t
Xbit_r115_c121 bl_121 br_121 wl_115 vdd gnd cell_6t
Xbit_r116_c121 bl_121 br_121 wl_116 vdd gnd cell_6t
Xbit_r117_c121 bl_121 br_121 wl_117 vdd gnd cell_6t
Xbit_r118_c121 bl_121 br_121 wl_118 vdd gnd cell_6t
Xbit_r119_c121 bl_121 br_121 wl_119 vdd gnd cell_6t
Xbit_r120_c121 bl_121 br_121 wl_120 vdd gnd cell_6t
Xbit_r121_c121 bl_121 br_121 wl_121 vdd gnd cell_6t
Xbit_r122_c121 bl_121 br_121 wl_122 vdd gnd cell_6t
Xbit_r123_c121 bl_121 br_121 wl_123 vdd gnd cell_6t
Xbit_r124_c121 bl_121 br_121 wl_124 vdd gnd cell_6t
Xbit_r125_c121 bl_121 br_121 wl_125 vdd gnd cell_6t
Xbit_r126_c121 bl_121 br_121 wl_126 vdd gnd cell_6t
Xbit_r127_c121 bl_121 br_121 wl_127 vdd gnd cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd cell_6t
Xbit_r1_c122 bl_122 br_122 wl_1 vdd gnd cell_6t
Xbit_r2_c122 bl_122 br_122 wl_2 vdd gnd cell_6t
Xbit_r3_c122 bl_122 br_122 wl_3 vdd gnd cell_6t
Xbit_r4_c122 bl_122 br_122 wl_4 vdd gnd cell_6t
Xbit_r5_c122 bl_122 br_122 wl_5 vdd gnd cell_6t
Xbit_r6_c122 bl_122 br_122 wl_6 vdd gnd cell_6t
Xbit_r7_c122 bl_122 br_122 wl_7 vdd gnd cell_6t
Xbit_r8_c122 bl_122 br_122 wl_8 vdd gnd cell_6t
Xbit_r9_c122 bl_122 br_122 wl_9 vdd gnd cell_6t
Xbit_r10_c122 bl_122 br_122 wl_10 vdd gnd cell_6t
Xbit_r11_c122 bl_122 br_122 wl_11 vdd gnd cell_6t
Xbit_r12_c122 bl_122 br_122 wl_12 vdd gnd cell_6t
Xbit_r13_c122 bl_122 br_122 wl_13 vdd gnd cell_6t
Xbit_r14_c122 bl_122 br_122 wl_14 vdd gnd cell_6t
Xbit_r15_c122 bl_122 br_122 wl_15 vdd gnd cell_6t
Xbit_r16_c122 bl_122 br_122 wl_16 vdd gnd cell_6t
Xbit_r17_c122 bl_122 br_122 wl_17 vdd gnd cell_6t
Xbit_r18_c122 bl_122 br_122 wl_18 vdd gnd cell_6t
Xbit_r19_c122 bl_122 br_122 wl_19 vdd gnd cell_6t
Xbit_r20_c122 bl_122 br_122 wl_20 vdd gnd cell_6t
Xbit_r21_c122 bl_122 br_122 wl_21 vdd gnd cell_6t
Xbit_r22_c122 bl_122 br_122 wl_22 vdd gnd cell_6t
Xbit_r23_c122 bl_122 br_122 wl_23 vdd gnd cell_6t
Xbit_r24_c122 bl_122 br_122 wl_24 vdd gnd cell_6t
Xbit_r25_c122 bl_122 br_122 wl_25 vdd gnd cell_6t
Xbit_r26_c122 bl_122 br_122 wl_26 vdd gnd cell_6t
Xbit_r27_c122 bl_122 br_122 wl_27 vdd gnd cell_6t
Xbit_r28_c122 bl_122 br_122 wl_28 vdd gnd cell_6t
Xbit_r29_c122 bl_122 br_122 wl_29 vdd gnd cell_6t
Xbit_r30_c122 bl_122 br_122 wl_30 vdd gnd cell_6t
Xbit_r31_c122 bl_122 br_122 wl_31 vdd gnd cell_6t
Xbit_r32_c122 bl_122 br_122 wl_32 vdd gnd cell_6t
Xbit_r33_c122 bl_122 br_122 wl_33 vdd gnd cell_6t
Xbit_r34_c122 bl_122 br_122 wl_34 vdd gnd cell_6t
Xbit_r35_c122 bl_122 br_122 wl_35 vdd gnd cell_6t
Xbit_r36_c122 bl_122 br_122 wl_36 vdd gnd cell_6t
Xbit_r37_c122 bl_122 br_122 wl_37 vdd gnd cell_6t
Xbit_r38_c122 bl_122 br_122 wl_38 vdd gnd cell_6t
Xbit_r39_c122 bl_122 br_122 wl_39 vdd gnd cell_6t
Xbit_r40_c122 bl_122 br_122 wl_40 vdd gnd cell_6t
Xbit_r41_c122 bl_122 br_122 wl_41 vdd gnd cell_6t
Xbit_r42_c122 bl_122 br_122 wl_42 vdd gnd cell_6t
Xbit_r43_c122 bl_122 br_122 wl_43 vdd gnd cell_6t
Xbit_r44_c122 bl_122 br_122 wl_44 vdd gnd cell_6t
Xbit_r45_c122 bl_122 br_122 wl_45 vdd gnd cell_6t
Xbit_r46_c122 bl_122 br_122 wl_46 vdd gnd cell_6t
Xbit_r47_c122 bl_122 br_122 wl_47 vdd gnd cell_6t
Xbit_r48_c122 bl_122 br_122 wl_48 vdd gnd cell_6t
Xbit_r49_c122 bl_122 br_122 wl_49 vdd gnd cell_6t
Xbit_r50_c122 bl_122 br_122 wl_50 vdd gnd cell_6t
Xbit_r51_c122 bl_122 br_122 wl_51 vdd gnd cell_6t
Xbit_r52_c122 bl_122 br_122 wl_52 vdd gnd cell_6t
Xbit_r53_c122 bl_122 br_122 wl_53 vdd gnd cell_6t
Xbit_r54_c122 bl_122 br_122 wl_54 vdd gnd cell_6t
Xbit_r55_c122 bl_122 br_122 wl_55 vdd gnd cell_6t
Xbit_r56_c122 bl_122 br_122 wl_56 vdd gnd cell_6t
Xbit_r57_c122 bl_122 br_122 wl_57 vdd gnd cell_6t
Xbit_r58_c122 bl_122 br_122 wl_58 vdd gnd cell_6t
Xbit_r59_c122 bl_122 br_122 wl_59 vdd gnd cell_6t
Xbit_r60_c122 bl_122 br_122 wl_60 vdd gnd cell_6t
Xbit_r61_c122 bl_122 br_122 wl_61 vdd gnd cell_6t
Xbit_r62_c122 bl_122 br_122 wl_62 vdd gnd cell_6t
Xbit_r63_c122 bl_122 br_122 wl_63 vdd gnd cell_6t
Xbit_r64_c122 bl_122 br_122 wl_64 vdd gnd cell_6t
Xbit_r65_c122 bl_122 br_122 wl_65 vdd gnd cell_6t
Xbit_r66_c122 bl_122 br_122 wl_66 vdd gnd cell_6t
Xbit_r67_c122 bl_122 br_122 wl_67 vdd gnd cell_6t
Xbit_r68_c122 bl_122 br_122 wl_68 vdd gnd cell_6t
Xbit_r69_c122 bl_122 br_122 wl_69 vdd gnd cell_6t
Xbit_r70_c122 bl_122 br_122 wl_70 vdd gnd cell_6t
Xbit_r71_c122 bl_122 br_122 wl_71 vdd gnd cell_6t
Xbit_r72_c122 bl_122 br_122 wl_72 vdd gnd cell_6t
Xbit_r73_c122 bl_122 br_122 wl_73 vdd gnd cell_6t
Xbit_r74_c122 bl_122 br_122 wl_74 vdd gnd cell_6t
Xbit_r75_c122 bl_122 br_122 wl_75 vdd gnd cell_6t
Xbit_r76_c122 bl_122 br_122 wl_76 vdd gnd cell_6t
Xbit_r77_c122 bl_122 br_122 wl_77 vdd gnd cell_6t
Xbit_r78_c122 bl_122 br_122 wl_78 vdd gnd cell_6t
Xbit_r79_c122 bl_122 br_122 wl_79 vdd gnd cell_6t
Xbit_r80_c122 bl_122 br_122 wl_80 vdd gnd cell_6t
Xbit_r81_c122 bl_122 br_122 wl_81 vdd gnd cell_6t
Xbit_r82_c122 bl_122 br_122 wl_82 vdd gnd cell_6t
Xbit_r83_c122 bl_122 br_122 wl_83 vdd gnd cell_6t
Xbit_r84_c122 bl_122 br_122 wl_84 vdd gnd cell_6t
Xbit_r85_c122 bl_122 br_122 wl_85 vdd gnd cell_6t
Xbit_r86_c122 bl_122 br_122 wl_86 vdd gnd cell_6t
Xbit_r87_c122 bl_122 br_122 wl_87 vdd gnd cell_6t
Xbit_r88_c122 bl_122 br_122 wl_88 vdd gnd cell_6t
Xbit_r89_c122 bl_122 br_122 wl_89 vdd gnd cell_6t
Xbit_r90_c122 bl_122 br_122 wl_90 vdd gnd cell_6t
Xbit_r91_c122 bl_122 br_122 wl_91 vdd gnd cell_6t
Xbit_r92_c122 bl_122 br_122 wl_92 vdd gnd cell_6t
Xbit_r93_c122 bl_122 br_122 wl_93 vdd gnd cell_6t
Xbit_r94_c122 bl_122 br_122 wl_94 vdd gnd cell_6t
Xbit_r95_c122 bl_122 br_122 wl_95 vdd gnd cell_6t
Xbit_r96_c122 bl_122 br_122 wl_96 vdd gnd cell_6t
Xbit_r97_c122 bl_122 br_122 wl_97 vdd gnd cell_6t
Xbit_r98_c122 bl_122 br_122 wl_98 vdd gnd cell_6t
Xbit_r99_c122 bl_122 br_122 wl_99 vdd gnd cell_6t
Xbit_r100_c122 bl_122 br_122 wl_100 vdd gnd cell_6t
Xbit_r101_c122 bl_122 br_122 wl_101 vdd gnd cell_6t
Xbit_r102_c122 bl_122 br_122 wl_102 vdd gnd cell_6t
Xbit_r103_c122 bl_122 br_122 wl_103 vdd gnd cell_6t
Xbit_r104_c122 bl_122 br_122 wl_104 vdd gnd cell_6t
Xbit_r105_c122 bl_122 br_122 wl_105 vdd gnd cell_6t
Xbit_r106_c122 bl_122 br_122 wl_106 vdd gnd cell_6t
Xbit_r107_c122 bl_122 br_122 wl_107 vdd gnd cell_6t
Xbit_r108_c122 bl_122 br_122 wl_108 vdd gnd cell_6t
Xbit_r109_c122 bl_122 br_122 wl_109 vdd gnd cell_6t
Xbit_r110_c122 bl_122 br_122 wl_110 vdd gnd cell_6t
Xbit_r111_c122 bl_122 br_122 wl_111 vdd gnd cell_6t
Xbit_r112_c122 bl_122 br_122 wl_112 vdd gnd cell_6t
Xbit_r113_c122 bl_122 br_122 wl_113 vdd gnd cell_6t
Xbit_r114_c122 bl_122 br_122 wl_114 vdd gnd cell_6t
Xbit_r115_c122 bl_122 br_122 wl_115 vdd gnd cell_6t
Xbit_r116_c122 bl_122 br_122 wl_116 vdd gnd cell_6t
Xbit_r117_c122 bl_122 br_122 wl_117 vdd gnd cell_6t
Xbit_r118_c122 bl_122 br_122 wl_118 vdd gnd cell_6t
Xbit_r119_c122 bl_122 br_122 wl_119 vdd gnd cell_6t
Xbit_r120_c122 bl_122 br_122 wl_120 vdd gnd cell_6t
Xbit_r121_c122 bl_122 br_122 wl_121 vdd gnd cell_6t
Xbit_r122_c122 bl_122 br_122 wl_122 vdd gnd cell_6t
Xbit_r123_c122 bl_122 br_122 wl_123 vdd gnd cell_6t
Xbit_r124_c122 bl_122 br_122 wl_124 vdd gnd cell_6t
Xbit_r125_c122 bl_122 br_122 wl_125 vdd gnd cell_6t
Xbit_r126_c122 bl_122 br_122 wl_126 vdd gnd cell_6t
Xbit_r127_c122 bl_122 br_122 wl_127 vdd gnd cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd cell_6t
Xbit_r1_c123 bl_123 br_123 wl_1 vdd gnd cell_6t
Xbit_r2_c123 bl_123 br_123 wl_2 vdd gnd cell_6t
Xbit_r3_c123 bl_123 br_123 wl_3 vdd gnd cell_6t
Xbit_r4_c123 bl_123 br_123 wl_4 vdd gnd cell_6t
Xbit_r5_c123 bl_123 br_123 wl_5 vdd gnd cell_6t
Xbit_r6_c123 bl_123 br_123 wl_6 vdd gnd cell_6t
Xbit_r7_c123 bl_123 br_123 wl_7 vdd gnd cell_6t
Xbit_r8_c123 bl_123 br_123 wl_8 vdd gnd cell_6t
Xbit_r9_c123 bl_123 br_123 wl_9 vdd gnd cell_6t
Xbit_r10_c123 bl_123 br_123 wl_10 vdd gnd cell_6t
Xbit_r11_c123 bl_123 br_123 wl_11 vdd gnd cell_6t
Xbit_r12_c123 bl_123 br_123 wl_12 vdd gnd cell_6t
Xbit_r13_c123 bl_123 br_123 wl_13 vdd gnd cell_6t
Xbit_r14_c123 bl_123 br_123 wl_14 vdd gnd cell_6t
Xbit_r15_c123 bl_123 br_123 wl_15 vdd gnd cell_6t
Xbit_r16_c123 bl_123 br_123 wl_16 vdd gnd cell_6t
Xbit_r17_c123 bl_123 br_123 wl_17 vdd gnd cell_6t
Xbit_r18_c123 bl_123 br_123 wl_18 vdd gnd cell_6t
Xbit_r19_c123 bl_123 br_123 wl_19 vdd gnd cell_6t
Xbit_r20_c123 bl_123 br_123 wl_20 vdd gnd cell_6t
Xbit_r21_c123 bl_123 br_123 wl_21 vdd gnd cell_6t
Xbit_r22_c123 bl_123 br_123 wl_22 vdd gnd cell_6t
Xbit_r23_c123 bl_123 br_123 wl_23 vdd gnd cell_6t
Xbit_r24_c123 bl_123 br_123 wl_24 vdd gnd cell_6t
Xbit_r25_c123 bl_123 br_123 wl_25 vdd gnd cell_6t
Xbit_r26_c123 bl_123 br_123 wl_26 vdd gnd cell_6t
Xbit_r27_c123 bl_123 br_123 wl_27 vdd gnd cell_6t
Xbit_r28_c123 bl_123 br_123 wl_28 vdd gnd cell_6t
Xbit_r29_c123 bl_123 br_123 wl_29 vdd gnd cell_6t
Xbit_r30_c123 bl_123 br_123 wl_30 vdd gnd cell_6t
Xbit_r31_c123 bl_123 br_123 wl_31 vdd gnd cell_6t
Xbit_r32_c123 bl_123 br_123 wl_32 vdd gnd cell_6t
Xbit_r33_c123 bl_123 br_123 wl_33 vdd gnd cell_6t
Xbit_r34_c123 bl_123 br_123 wl_34 vdd gnd cell_6t
Xbit_r35_c123 bl_123 br_123 wl_35 vdd gnd cell_6t
Xbit_r36_c123 bl_123 br_123 wl_36 vdd gnd cell_6t
Xbit_r37_c123 bl_123 br_123 wl_37 vdd gnd cell_6t
Xbit_r38_c123 bl_123 br_123 wl_38 vdd gnd cell_6t
Xbit_r39_c123 bl_123 br_123 wl_39 vdd gnd cell_6t
Xbit_r40_c123 bl_123 br_123 wl_40 vdd gnd cell_6t
Xbit_r41_c123 bl_123 br_123 wl_41 vdd gnd cell_6t
Xbit_r42_c123 bl_123 br_123 wl_42 vdd gnd cell_6t
Xbit_r43_c123 bl_123 br_123 wl_43 vdd gnd cell_6t
Xbit_r44_c123 bl_123 br_123 wl_44 vdd gnd cell_6t
Xbit_r45_c123 bl_123 br_123 wl_45 vdd gnd cell_6t
Xbit_r46_c123 bl_123 br_123 wl_46 vdd gnd cell_6t
Xbit_r47_c123 bl_123 br_123 wl_47 vdd gnd cell_6t
Xbit_r48_c123 bl_123 br_123 wl_48 vdd gnd cell_6t
Xbit_r49_c123 bl_123 br_123 wl_49 vdd gnd cell_6t
Xbit_r50_c123 bl_123 br_123 wl_50 vdd gnd cell_6t
Xbit_r51_c123 bl_123 br_123 wl_51 vdd gnd cell_6t
Xbit_r52_c123 bl_123 br_123 wl_52 vdd gnd cell_6t
Xbit_r53_c123 bl_123 br_123 wl_53 vdd gnd cell_6t
Xbit_r54_c123 bl_123 br_123 wl_54 vdd gnd cell_6t
Xbit_r55_c123 bl_123 br_123 wl_55 vdd gnd cell_6t
Xbit_r56_c123 bl_123 br_123 wl_56 vdd gnd cell_6t
Xbit_r57_c123 bl_123 br_123 wl_57 vdd gnd cell_6t
Xbit_r58_c123 bl_123 br_123 wl_58 vdd gnd cell_6t
Xbit_r59_c123 bl_123 br_123 wl_59 vdd gnd cell_6t
Xbit_r60_c123 bl_123 br_123 wl_60 vdd gnd cell_6t
Xbit_r61_c123 bl_123 br_123 wl_61 vdd gnd cell_6t
Xbit_r62_c123 bl_123 br_123 wl_62 vdd gnd cell_6t
Xbit_r63_c123 bl_123 br_123 wl_63 vdd gnd cell_6t
Xbit_r64_c123 bl_123 br_123 wl_64 vdd gnd cell_6t
Xbit_r65_c123 bl_123 br_123 wl_65 vdd gnd cell_6t
Xbit_r66_c123 bl_123 br_123 wl_66 vdd gnd cell_6t
Xbit_r67_c123 bl_123 br_123 wl_67 vdd gnd cell_6t
Xbit_r68_c123 bl_123 br_123 wl_68 vdd gnd cell_6t
Xbit_r69_c123 bl_123 br_123 wl_69 vdd gnd cell_6t
Xbit_r70_c123 bl_123 br_123 wl_70 vdd gnd cell_6t
Xbit_r71_c123 bl_123 br_123 wl_71 vdd gnd cell_6t
Xbit_r72_c123 bl_123 br_123 wl_72 vdd gnd cell_6t
Xbit_r73_c123 bl_123 br_123 wl_73 vdd gnd cell_6t
Xbit_r74_c123 bl_123 br_123 wl_74 vdd gnd cell_6t
Xbit_r75_c123 bl_123 br_123 wl_75 vdd gnd cell_6t
Xbit_r76_c123 bl_123 br_123 wl_76 vdd gnd cell_6t
Xbit_r77_c123 bl_123 br_123 wl_77 vdd gnd cell_6t
Xbit_r78_c123 bl_123 br_123 wl_78 vdd gnd cell_6t
Xbit_r79_c123 bl_123 br_123 wl_79 vdd gnd cell_6t
Xbit_r80_c123 bl_123 br_123 wl_80 vdd gnd cell_6t
Xbit_r81_c123 bl_123 br_123 wl_81 vdd gnd cell_6t
Xbit_r82_c123 bl_123 br_123 wl_82 vdd gnd cell_6t
Xbit_r83_c123 bl_123 br_123 wl_83 vdd gnd cell_6t
Xbit_r84_c123 bl_123 br_123 wl_84 vdd gnd cell_6t
Xbit_r85_c123 bl_123 br_123 wl_85 vdd gnd cell_6t
Xbit_r86_c123 bl_123 br_123 wl_86 vdd gnd cell_6t
Xbit_r87_c123 bl_123 br_123 wl_87 vdd gnd cell_6t
Xbit_r88_c123 bl_123 br_123 wl_88 vdd gnd cell_6t
Xbit_r89_c123 bl_123 br_123 wl_89 vdd gnd cell_6t
Xbit_r90_c123 bl_123 br_123 wl_90 vdd gnd cell_6t
Xbit_r91_c123 bl_123 br_123 wl_91 vdd gnd cell_6t
Xbit_r92_c123 bl_123 br_123 wl_92 vdd gnd cell_6t
Xbit_r93_c123 bl_123 br_123 wl_93 vdd gnd cell_6t
Xbit_r94_c123 bl_123 br_123 wl_94 vdd gnd cell_6t
Xbit_r95_c123 bl_123 br_123 wl_95 vdd gnd cell_6t
Xbit_r96_c123 bl_123 br_123 wl_96 vdd gnd cell_6t
Xbit_r97_c123 bl_123 br_123 wl_97 vdd gnd cell_6t
Xbit_r98_c123 bl_123 br_123 wl_98 vdd gnd cell_6t
Xbit_r99_c123 bl_123 br_123 wl_99 vdd gnd cell_6t
Xbit_r100_c123 bl_123 br_123 wl_100 vdd gnd cell_6t
Xbit_r101_c123 bl_123 br_123 wl_101 vdd gnd cell_6t
Xbit_r102_c123 bl_123 br_123 wl_102 vdd gnd cell_6t
Xbit_r103_c123 bl_123 br_123 wl_103 vdd gnd cell_6t
Xbit_r104_c123 bl_123 br_123 wl_104 vdd gnd cell_6t
Xbit_r105_c123 bl_123 br_123 wl_105 vdd gnd cell_6t
Xbit_r106_c123 bl_123 br_123 wl_106 vdd gnd cell_6t
Xbit_r107_c123 bl_123 br_123 wl_107 vdd gnd cell_6t
Xbit_r108_c123 bl_123 br_123 wl_108 vdd gnd cell_6t
Xbit_r109_c123 bl_123 br_123 wl_109 vdd gnd cell_6t
Xbit_r110_c123 bl_123 br_123 wl_110 vdd gnd cell_6t
Xbit_r111_c123 bl_123 br_123 wl_111 vdd gnd cell_6t
Xbit_r112_c123 bl_123 br_123 wl_112 vdd gnd cell_6t
Xbit_r113_c123 bl_123 br_123 wl_113 vdd gnd cell_6t
Xbit_r114_c123 bl_123 br_123 wl_114 vdd gnd cell_6t
Xbit_r115_c123 bl_123 br_123 wl_115 vdd gnd cell_6t
Xbit_r116_c123 bl_123 br_123 wl_116 vdd gnd cell_6t
Xbit_r117_c123 bl_123 br_123 wl_117 vdd gnd cell_6t
Xbit_r118_c123 bl_123 br_123 wl_118 vdd gnd cell_6t
Xbit_r119_c123 bl_123 br_123 wl_119 vdd gnd cell_6t
Xbit_r120_c123 bl_123 br_123 wl_120 vdd gnd cell_6t
Xbit_r121_c123 bl_123 br_123 wl_121 vdd gnd cell_6t
Xbit_r122_c123 bl_123 br_123 wl_122 vdd gnd cell_6t
Xbit_r123_c123 bl_123 br_123 wl_123 vdd gnd cell_6t
Xbit_r124_c123 bl_123 br_123 wl_124 vdd gnd cell_6t
Xbit_r125_c123 bl_123 br_123 wl_125 vdd gnd cell_6t
Xbit_r126_c123 bl_123 br_123 wl_126 vdd gnd cell_6t
Xbit_r127_c123 bl_123 br_123 wl_127 vdd gnd cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd cell_6t
Xbit_r1_c124 bl_124 br_124 wl_1 vdd gnd cell_6t
Xbit_r2_c124 bl_124 br_124 wl_2 vdd gnd cell_6t
Xbit_r3_c124 bl_124 br_124 wl_3 vdd gnd cell_6t
Xbit_r4_c124 bl_124 br_124 wl_4 vdd gnd cell_6t
Xbit_r5_c124 bl_124 br_124 wl_5 vdd gnd cell_6t
Xbit_r6_c124 bl_124 br_124 wl_6 vdd gnd cell_6t
Xbit_r7_c124 bl_124 br_124 wl_7 vdd gnd cell_6t
Xbit_r8_c124 bl_124 br_124 wl_8 vdd gnd cell_6t
Xbit_r9_c124 bl_124 br_124 wl_9 vdd gnd cell_6t
Xbit_r10_c124 bl_124 br_124 wl_10 vdd gnd cell_6t
Xbit_r11_c124 bl_124 br_124 wl_11 vdd gnd cell_6t
Xbit_r12_c124 bl_124 br_124 wl_12 vdd gnd cell_6t
Xbit_r13_c124 bl_124 br_124 wl_13 vdd gnd cell_6t
Xbit_r14_c124 bl_124 br_124 wl_14 vdd gnd cell_6t
Xbit_r15_c124 bl_124 br_124 wl_15 vdd gnd cell_6t
Xbit_r16_c124 bl_124 br_124 wl_16 vdd gnd cell_6t
Xbit_r17_c124 bl_124 br_124 wl_17 vdd gnd cell_6t
Xbit_r18_c124 bl_124 br_124 wl_18 vdd gnd cell_6t
Xbit_r19_c124 bl_124 br_124 wl_19 vdd gnd cell_6t
Xbit_r20_c124 bl_124 br_124 wl_20 vdd gnd cell_6t
Xbit_r21_c124 bl_124 br_124 wl_21 vdd gnd cell_6t
Xbit_r22_c124 bl_124 br_124 wl_22 vdd gnd cell_6t
Xbit_r23_c124 bl_124 br_124 wl_23 vdd gnd cell_6t
Xbit_r24_c124 bl_124 br_124 wl_24 vdd gnd cell_6t
Xbit_r25_c124 bl_124 br_124 wl_25 vdd gnd cell_6t
Xbit_r26_c124 bl_124 br_124 wl_26 vdd gnd cell_6t
Xbit_r27_c124 bl_124 br_124 wl_27 vdd gnd cell_6t
Xbit_r28_c124 bl_124 br_124 wl_28 vdd gnd cell_6t
Xbit_r29_c124 bl_124 br_124 wl_29 vdd gnd cell_6t
Xbit_r30_c124 bl_124 br_124 wl_30 vdd gnd cell_6t
Xbit_r31_c124 bl_124 br_124 wl_31 vdd gnd cell_6t
Xbit_r32_c124 bl_124 br_124 wl_32 vdd gnd cell_6t
Xbit_r33_c124 bl_124 br_124 wl_33 vdd gnd cell_6t
Xbit_r34_c124 bl_124 br_124 wl_34 vdd gnd cell_6t
Xbit_r35_c124 bl_124 br_124 wl_35 vdd gnd cell_6t
Xbit_r36_c124 bl_124 br_124 wl_36 vdd gnd cell_6t
Xbit_r37_c124 bl_124 br_124 wl_37 vdd gnd cell_6t
Xbit_r38_c124 bl_124 br_124 wl_38 vdd gnd cell_6t
Xbit_r39_c124 bl_124 br_124 wl_39 vdd gnd cell_6t
Xbit_r40_c124 bl_124 br_124 wl_40 vdd gnd cell_6t
Xbit_r41_c124 bl_124 br_124 wl_41 vdd gnd cell_6t
Xbit_r42_c124 bl_124 br_124 wl_42 vdd gnd cell_6t
Xbit_r43_c124 bl_124 br_124 wl_43 vdd gnd cell_6t
Xbit_r44_c124 bl_124 br_124 wl_44 vdd gnd cell_6t
Xbit_r45_c124 bl_124 br_124 wl_45 vdd gnd cell_6t
Xbit_r46_c124 bl_124 br_124 wl_46 vdd gnd cell_6t
Xbit_r47_c124 bl_124 br_124 wl_47 vdd gnd cell_6t
Xbit_r48_c124 bl_124 br_124 wl_48 vdd gnd cell_6t
Xbit_r49_c124 bl_124 br_124 wl_49 vdd gnd cell_6t
Xbit_r50_c124 bl_124 br_124 wl_50 vdd gnd cell_6t
Xbit_r51_c124 bl_124 br_124 wl_51 vdd gnd cell_6t
Xbit_r52_c124 bl_124 br_124 wl_52 vdd gnd cell_6t
Xbit_r53_c124 bl_124 br_124 wl_53 vdd gnd cell_6t
Xbit_r54_c124 bl_124 br_124 wl_54 vdd gnd cell_6t
Xbit_r55_c124 bl_124 br_124 wl_55 vdd gnd cell_6t
Xbit_r56_c124 bl_124 br_124 wl_56 vdd gnd cell_6t
Xbit_r57_c124 bl_124 br_124 wl_57 vdd gnd cell_6t
Xbit_r58_c124 bl_124 br_124 wl_58 vdd gnd cell_6t
Xbit_r59_c124 bl_124 br_124 wl_59 vdd gnd cell_6t
Xbit_r60_c124 bl_124 br_124 wl_60 vdd gnd cell_6t
Xbit_r61_c124 bl_124 br_124 wl_61 vdd gnd cell_6t
Xbit_r62_c124 bl_124 br_124 wl_62 vdd gnd cell_6t
Xbit_r63_c124 bl_124 br_124 wl_63 vdd gnd cell_6t
Xbit_r64_c124 bl_124 br_124 wl_64 vdd gnd cell_6t
Xbit_r65_c124 bl_124 br_124 wl_65 vdd gnd cell_6t
Xbit_r66_c124 bl_124 br_124 wl_66 vdd gnd cell_6t
Xbit_r67_c124 bl_124 br_124 wl_67 vdd gnd cell_6t
Xbit_r68_c124 bl_124 br_124 wl_68 vdd gnd cell_6t
Xbit_r69_c124 bl_124 br_124 wl_69 vdd gnd cell_6t
Xbit_r70_c124 bl_124 br_124 wl_70 vdd gnd cell_6t
Xbit_r71_c124 bl_124 br_124 wl_71 vdd gnd cell_6t
Xbit_r72_c124 bl_124 br_124 wl_72 vdd gnd cell_6t
Xbit_r73_c124 bl_124 br_124 wl_73 vdd gnd cell_6t
Xbit_r74_c124 bl_124 br_124 wl_74 vdd gnd cell_6t
Xbit_r75_c124 bl_124 br_124 wl_75 vdd gnd cell_6t
Xbit_r76_c124 bl_124 br_124 wl_76 vdd gnd cell_6t
Xbit_r77_c124 bl_124 br_124 wl_77 vdd gnd cell_6t
Xbit_r78_c124 bl_124 br_124 wl_78 vdd gnd cell_6t
Xbit_r79_c124 bl_124 br_124 wl_79 vdd gnd cell_6t
Xbit_r80_c124 bl_124 br_124 wl_80 vdd gnd cell_6t
Xbit_r81_c124 bl_124 br_124 wl_81 vdd gnd cell_6t
Xbit_r82_c124 bl_124 br_124 wl_82 vdd gnd cell_6t
Xbit_r83_c124 bl_124 br_124 wl_83 vdd gnd cell_6t
Xbit_r84_c124 bl_124 br_124 wl_84 vdd gnd cell_6t
Xbit_r85_c124 bl_124 br_124 wl_85 vdd gnd cell_6t
Xbit_r86_c124 bl_124 br_124 wl_86 vdd gnd cell_6t
Xbit_r87_c124 bl_124 br_124 wl_87 vdd gnd cell_6t
Xbit_r88_c124 bl_124 br_124 wl_88 vdd gnd cell_6t
Xbit_r89_c124 bl_124 br_124 wl_89 vdd gnd cell_6t
Xbit_r90_c124 bl_124 br_124 wl_90 vdd gnd cell_6t
Xbit_r91_c124 bl_124 br_124 wl_91 vdd gnd cell_6t
Xbit_r92_c124 bl_124 br_124 wl_92 vdd gnd cell_6t
Xbit_r93_c124 bl_124 br_124 wl_93 vdd gnd cell_6t
Xbit_r94_c124 bl_124 br_124 wl_94 vdd gnd cell_6t
Xbit_r95_c124 bl_124 br_124 wl_95 vdd gnd cell_6t
Xbit_r96_c124 bl_124 br_124 wl_96 vdd gnd cell_6t
Xbit_r97_c124 bl_124 br_124 wl_97 vdd gnd cell_6t
Xbit_r98_c124 bl_124 br_124 wl_98 vdd gnd cell_6t
Xbit_r99_c124 bl_124 br_124 wl_99 vdd gnd cell_6t
Xbit_r100_c124 bl_124 br_124 wl_100 vdd gnd cell_6t
Xbit_r101_c124 bl_124 br_124 wl_101 vdd gnd cell_6t
Xbit_r102_c124 bl_124 br_124 wl_102 vdd gnd cell_6t
Xbit_r103_c124 bl_124 br_124 wl_103 vdd gnd cell_6t
Xbit_r104_c124 bl_124 br_124 wl_104 vdd gnd cell_6t
Xbit_r105_c124 bl_124 br_124 wl_105 vdd gnd cell_6t
Xbit_r106_c124 bl_124 br_124 wl_106 vdd gnd cell_6t
Xbit_r107_c124 bl_124 br_124 wl_107 vdd gnd cell_6t
Xbit_r108_c124 bl_124 br_124 wl_108 vdd gnd cell_6t
Xbit_r109_c124 bl_124 br_124 wl_109 vdd gnd cell_6t
Xbit_r110_c124 bl_124 br_124 wl_110 vdd gnd cell_6t
Xbit_r111_c124 bl_124 br_124 wl_111 vdd gnd cell_6t
Xbit_r112_c124 bl_124 br_124 wl_112 vdd gnd cell_6t
Xbit_r113_c124 bl_124 br_124 wl_113 vdd gnd cell_6t
Xbit_r114_c124 bl_124 br_124 wl_114 vdd gnd cell_6t
Xbit_r115_c124 bl_124 br_124 wl_115 vdd gnd cell_6t
Xbit_r116_c124 bl_124 br_124 wl_116 vdd gnd cell_6t
Xbit_r117_c124 bl_124 br_124 wl_117 vdd gnd cell_6t
Xbit_r118_c124 bl_124 br_124 wl_118 vdd gnd cell_6t
Xbit_r119_c124 bl_124 br_124 wl_119 vdd gnd cell_6t
Xbit_r120_c124 bl_124 br_124 wl_120 vdd gnd cell_6t
Xbit_r121_c124 bl_124 br_124 wl_121 vdd gnd cell_6t
Xbit_r122_c124 bl_124 br_124 wl_122 vdd gnd cell_6t
Xbit_r123_c124 bl_124 br_124 wl_123 vdd gnd cell_6t
Xbit_r124_c124 bl_124 br_124 wl_124 vdd gnd cell_6t
Xbit_r125_c124 bl_124 br_124 wl_125 vdd gnd cell_6t
Xbit_r126_c124 bl_124 br_124 wl_126 vdd gnd cell_6t
Xbit_r127_c124 bl_124 br_124 wl_127 vdd gnd cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd cell_6t
Xbit_r1_c125 bl_125 br_125 wl_1 vdd gnd cell_6t
Xbit_r2_c125 bl_125 br_125 wl_2 vdd gnd cell_6t
Xbit_r3_c125 bl_125 br_125 wl_3 vdd gnd cell_6t
Xbit_r4_c125 bl_125 br_125 wl_4 vdd gnd cell_6t
Xbit_r5_c125 bl_125 br_125 wl_5 vdd gnd cell_6t
Xbit_r6_c125 bl_125 br_125 wl_6 vdd gnd cell_6t
Xbit_r7_c125 bl_125 br_125 wl_7 vdd gnd cell_6t
Xbit_r8_c125 bl_125 br_125 wl_8 vdd gnd cell_6t
Xbit_r9_c125 bl_125 br_125 wl_9 vdd gnd cell_6t
Xbit_r10_c125 bl_125 br_125 wl_10 vdd gnd cell_6t
Xbit_r11_c125 bl_125 br_125 wl_11 vdd gnd cell_6t
Xbit_r12_c125 bl_125 br_125 wl_12 vdd gnd cell_6t
Xbit_r13_c125 bl_125 br_125 wl_13 vdd gnd cell_6t
Xbit_r14_c125 bl_125 br_125 wl_14 vdd gnd cell_6t
Xbit_r15_c125 bl_125 br_125 wl_15 vdd gnd cell_6t
Xbit_r16_c125 bl_125 br_125 wl_16 vdd gnd cell_6t
Xbit_r17_c125 bl_125 br_125 wl_17 vdd gnd cell_6t
Xbit_r18_c125 bl_125 br_125 wl_18 vdd gnd cell_6t
Xbit_r19_c125 bl_125 br_125 wl_19 vdd gnd cell_6t
Xbit_r20_c125 bl_125 br_125 wl_20 vdd gnd cell_6t
Xbit_r21_c125 bl_125 br_125 wl_21 vdd gnd cell_6t
Xbit_r22_c125 bl_125 br_125 wl_22 vdd gnd cell_6t
Xbit_r23_c125 bl_125 br_125 wl_23 vdd gnd cell_6t
Xbit_r24_c125 bl_125 br_125 wl_24 vdd gnd cell_6t
Xbit_r25_c125 bl_125 br_125 wl_25 vdd gnd cell_6t
Xbit_r26_c125 bl_125 br_125 wl_26 vdd gnd cell_6t
Xbit_r27_c125 bl_125 br_125 wl_27 vdd gnd cell_6t
Xbit_r28_c125 bl_125 br_125 wl_28 vdd gnd cell_6t
Xbit_r29_c125 bl_125 br_125 wl_29 vdd gnd cell_6t
Xbit_r30_c125 bl_125 br_125 wl_30 vdd gnd cell_6t
Xbit_r31_c125 bl_125 br_125 wl_31 vdd gnd cell_6t
Xbit_r32_c125 bl_125 br_125 wl_32 vdd gnd cell_6t
Xbit_r33_c125 bl_125 br_125 wl_33 vdd gnd cell_6t
Xbit_r34_c125 bl_125 br_125 wl_34 vdd gnd cell_6t
Xbit_r35_c125 bl_125 br_125 wl_35 vdd gnd cell_6t
Xbit_r36_c125 bl_125 br_125 wl_36 vdd gnd cell_6t
Xbit_r37_c125 bl_125 br_125 wl_37 vdd gnd cell_6t
Xbit_r38_c125 bl_125 br_125 wl_38 vdd gnd cell_6t
Xbit_r39_c125 bl_125 br_125 wl_39 vdd gnd cell_6t
Xbit_r40_c125 bl_125 br_125 wl_40 vdd gnd cell_6t
Xbit_r41_c125 bl_125 br_125 wl_41 vdd gnd cell_6t
Xbit_r42_c125 bl_125 br_125 wl_42 vdd gnd cell_6t
Xbit_r43_c125 bl_125 br_125 wl_43 vdd gnd cell_6t
Xbit_r44_c125 bl_125 br_125 wl_44 vdd gnd cell_6t
Xbit_r45_c125 bl_125 br_125 wl_45 vdd gnd cell_6t
Xbit_r46_c125 bl_125 br_125 wl_46 vdd gnd cell_6t
Xbit_r47_c125 bl_125 br_125 wl_47 vdd gnd cell_6t
Xbit_r48_c125 bl_125 br_125 wl_48 vdd gnd cell_6t
Xbit_r49_c125 bl_125 br_125 wl_49 vdd gnd cell_6t
Xbit_r50_c125 bl_125 br_125 wl_50 vdd gnd cell_6t
Xbit_r51_c125 bl_125 br_125 wl_51 vdd gnd cell_6t
Xbit_r52_c125 bl_125 br_125 wl_52 vdd gnd cell_6t
Xbit_r53_c125 bl_125 br_125 wl_53 vdd gnd cell_6t
Xbit_r54_c125 bl_125 br_125 wl_54 vdd gnd cell_6t
Xbit_r55_c125 bl_125 br_125 wl_55 vdd gnd cell_6t
Xbit_r56_c125 bl_125 br_125 wl_56 vdd gnd cell_6t
Xbit_r57_c125 bl_125 br_125 wl_57 vdd gnd cell_6t
Xbit_r58_c125 bl_125 br_125 wl_58 vdd gnd cell_6t
Xbit_r59_c125 bl_125 br_125 wl_59 vdd gnd cell_6t
Xbit_r60_c125 bl_125 br_125 wl_60 vdd gnd cell_6t
Xbit_r61_c125 bl_125 br_125 wl_61 vdd gnd cell_6t
Xbit_r62_c125 bl_125 br_125 wl_62 vdd gnd cell_6t
Xbit_r63_c125 bl_125 br_125 wl_63 vdd gnd cell_6t
Xbit_r64_c125 bl_125 br_125 wl_64 vdd gnd cell_6t
Xbit_r65_c125 bl_125 br_125 wl_65 vdd gnd cell_6t
Xbit_r66_c125 bl_125 br_125 wl_66 vdd gnd cell_6t
Xbit_r67_c125 bl_125 br_125 wl_67 vdd gnd cell_6t
Xbit_r68_c125 bl_125 br_125 wl_68 vdd gnd cell_6t
Xbit_r69_c125 bl_125 br_125 wl_69 vdd gnd cell_6t
Xbit_r70_c125 bl_125 br_125 wl_70 vdd gnd cell_6t
Xbit_r71_c125 bl_125 br_125 wl_71 vdd gnd cell_6t
Xbit_r72_c125 bl_125 br_125 wl_72 vdd gnd cell_6t
Xbit_r73_c125 bl_125 br_125 wl_73 vdd gnd cell_6t
Xbit_r74_c125 bl_125 br_125 wl_74 vdd gnd cell_6t
Xbit_r75_c125 bl_125 br_125 wl_75 vdd gnd cell_6t
Xbit_r76_c125 bl_125 br_125 wl_76 vdd gnd cell_6t
Xbit_r77_c125 bl_125 br_125 wl_77 vdd gnd cell_6t
Xbit_r78_c125 bl_125 br_125 wl_78 vdd gnd cell_6t
Xbit_r79_c125 bl_125 br_125 wl_79 vdd gnd cell_6t
Xbit_r80_c125 bl_125 br_125 wl_80 vdd gnd cell_6t
Xbit_r81_c125 bl_125 br_125 wl_81 vdd gnd cell_6t
Xbit_r82_c125 bl_125 br_125 wl_82 vdd gnd cell_6t
Xbit_r83_c125 bl_125 br_125 wl_83 vdd gnd cell_6t
Xbit_r84_c125 bl_125 br_125 wl_84 vdd gnd cell_6t
Xbit_r85_c125 bl_125 br_125 wl_85 vdd gnd cell_6t
Xbit_r86_c125 bl_125 br_125 wl_86 vdd gnd cell_6t
Xbit_r87_c125 bl_125 br_125 wl_87 vdd gnd cell_6t
Xbit_r88_c125 bl_125 br_125 wl_88 vdd gnd cell_6t
Xbit_r89_c125 bl_125 br_125 wl_89 vdd gnd cell_6t
Xbit_r90_c125 bl_125 br_125 wl_90 vdd gnd cell_6t
Xbit_r91_c125 bl_125 br_125 wl_91 vdd gnd cell_6t
Xbit_r92_c125 bl_125 br_125 wl_92 vdd gnd cell_6t
Xbit_r93_c125 bl_125 br_125 wl_93 vdd gnd cell_6t
Xbit_r94_c125 bl_125 br_125 wl_94 vdd gnd cell_6t
Xbit_r95_c125 bl_125 br_125 wl_95 vdd gnd cell_6t
Xbit_r96_c125 bl_125 br_125 wl_96 vdd gnd cell_6t
Xbit_r97_c125 bl_125 br_125 wl_97 vdd gnd cell_6t
Xbit_r98_c125 bl_125 br_125 wl_98 vdd gnd cell_6t
Xbit_r99_c125 bl_125 br_125 wl_99 vdd gnd cell_6t
Xbit_r100_c125 bl_125 br_125 wl_100 vdd gnd cell_6t
Xbit_r101_c125 bl_125 br_125 wl_101 vdd gnd cell_6t
Xbit_r102_c125 bl_125 br_125 wl_102 vdd gnd cell_6t
Xbit_r103_c125 bl_125 br_125 wl_103 vdd gnd cell_6t
Xbit_r104_c125 bl_125 br_125 wl_104 vdd gnd cell_6t
Xbit_r105_c125 bl_125 br_125 wl_105 vdd gnd cell_6t
Xbit_r106_c125 bl_125 br_125 wl_106 vdd gnd cell_6t
Xbit_r107_c125 bl_125 br_125 wl_107 vdd gnd cell_6t
Xbit_r108_c125 bl_125 br_125 wl_108 vdd gnd cell_6t
Xbit_r109_c125 bl_125 br_125 wl_109 vdd gnd cell_6t
Xbit_r110_c125 bl_125 br_125 wl_110 vdd gnd cell_6t
Xbit_r111_c125 bl_125 br_125 wl_111 vdd gnd cell_6t
Xbit_r112_c125 bl_125 br_125 wl_112 vdd gnd cell_6t
Xbit_r113_c125 bl_125 br_125 wl_113 vdd gnd cell_6t
Xbit_r114_c125 bl_125 br_125 wl_114 vdd gnd cell_6t
Xbit_r115_c125 bl_125 br_125 wl_115 vdd gnd cell_6t
Xbit_r116_c125 bl_125 br_125 wl_116 vdd gnd cell_6t
Xbit_r117_c125 bl_125 br_125 wl_117 vdd gnd cell_6t
Xbit_r118_c125 bl_125 br_125 wl_118 vdd gnd cell_6t
Xbit_r119_c125 bl_125 br_125 wl_119 vdd gnd cell_6t
Xbit_r120_c125 bl_125 br_125 wl_120 vdd gnd cell_6t
Xbit_r121_c125 bl_125 br_125 wl_121 vdd gnd cell_6t
Xbit_r122_c125 bl_125 br_125 wl_122 vdd gnd cell_6t
Xbit_r123_c125 bl_125 br_125 wl_123 vdd gnd cell_6t
Xbit_r124_c125 bl_125 br_125 wl_124 vdd gnd cell_6t
Xbit_r125_c125 bl_125 br_125 wl_125 vdd gnd cell_6t
Xbit_r126_c125 bl_125 br_125 wl_126 vdd gnd cell_6t
Xbit_r127_c125 bl_125 br_125 wl_127 vdd gnd cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd cell_6t
Xbit_r1_c126 bl_126 br_126 wl_1 vdd gnd cell_6t
Xbit_r2_c126 bl_126 br_126 wl_2 vdd gnd cell_6t
Xbit_r3_c126 bl_126 br_126 wl_3 vdd gnd cell_6t
Xbit_r4_c126 bl_126 br_126 wl_4 vdd gnd cell_6t
Xbit_r5_c126 bl_126 br_126 wl_5 vdd gnd cell_6t
Xbit_r6_c126 bl_126 br_126 wl_6 vdd gnd cell_6t
Xbit_r7_c126 bl_126 br_126 wl_7 vdd gnd cell_6t
Xbit_r8_c126 bl_126 br_126 wl_8 vdd gnd cell_6t
Xbit_r9_c126 bl_126 br_126 wl_9 vdd gnd cell_6t
Xbit_r10_c126 bl_126 br_126 wl_10 vdd gnd cell_6t
Xbit_r11_c126 bl_126 br_126 wl_11 vdd gnd cell_6t
Xbit_r12_c126 bl_126 br_126 wl_12 vdd gnd cell_6t
Xbit_r13_c126 bl_126 br_126 wl_13 vdd gnd cell_6t
Xbit_r14_c126 bl_126 br_126 wl_14 vdd gnd cell_6t
Xbit_r15_c126 bl_126 br_126 wl_15 vdd gnd cell_6t
Xbit_r16_c126 bl_126 br_126 wl_16 vdd gnd cell_6t
Xbit_r17_c126 bl_126 br_126 wl_17 vdd gnd cell_6t
Xbit_r18_c126 bl_126 br_126 wl_18 vdd gnd cell_6t
Xbit_r19_c126 bl_126 br_126 wl_19 vdd gnd cell_6t
Xbit_r20_c126 bl_126 br_126 wl_20 vdd gnd cell_6t
Xbit_r21_c126 bl_126 br_126 wl_21 vdd gnd cell_6t
Xbit_r22_c126 bl_126 br_126 wl_22 vdd gnd cell_6t
Xbit_r23_c126 bl_126 br_126 wl_23 vdd gnd cell_6t
Xbit_r24_c126 bl_126 br_126 wl_24 vdd gnd cell_6t
Xbit_r25_c126 bl_126 br_126 wl_25 vdd gnd cell_6t
Xbit_r26_c126 bl_126 br_126 wl_26 vdd gnd cell_6t
Xbit_r27_c126 bl_126 br_126 wl_27 vdd gnd cell_6t
Xbit_r28_c126 bl_126 br_126 wl_28 vdd gnd cell_6t
Xbit_r29_c126 bl_126 br_126 wl_29 vdd gnd cell_6t
Xbit_r30_c126 bl_126 br_126 wl_30 vdd gnd cell_6t
Xbit_r31_c126 bl_126 br_126 wl_31 vdd gnd cell_6t
Xbit_r32_c126 bl_126 br_126 wl_32 vdd gnd cell_6t
Xbit_r33_c126 bl_126 br_126 wl_33 vdd gnd cell_6t
Xbit_r34_c126 bl_126 br_126 wl_34 vdd gnd cell_6t
Xbit_r35_c126 bl_126 br_126 wl_35 vdd gnd cell_6t
Xbit_r36_c126 bl_126 br_126 wl_36 vdd gnd cell_6t
Xbit_r37_c126 bl_126 br_126 wl_37 vdd gnd cell_6t
Xbit_r38_c126 bl_126 br_126 wl_38 vdd gnd cell_6t
Xbit_r39_c126 bl_126 br_126 wl_39 vdd gnd cell_6t
Xbit_r40_c126 bl_126 br_126 wl_40 vdd gnd cell_6t
Xbit_r41_c126 bl_126 br_126 wl_41 vdd gnd cell_6t
Xbit_r42_c126 bl_126 br_126 wl_42 vdd gnd cell_6t
Xbit_r43_c126 bl_126 br_126 wl_43 vdd gnd cell_6t
Xbit_r44_c126 bl_126 br_126 wl_44 vdd gnd cell_6t
Xbit_r45_c126 bl_126 br_126 wl_45 vdd gnd cell_6t
Xbit_r46_c126 bl_126 br_126 wl_46 vdd gnd cell_6t
Xbit_r47_c126 bl_126 br_126 wl_47 vdd gnd cell_6t
Xbit_r48_c126 bl_126 br_126 wl_48 vdd gnd cell_6t
Xbit_r49_c126 bl_126 br_126 wl_49 vdd gnd cell_6t
Xbit_r50_c126 bl_126 br_126 wl_50 vdd gnd cell_6t
Xbit_r51_c126 bl_126 br_126 wl_51 vdd gnd cell_6t
Xbit_r52_c126 bl_126 br_126 wl_52 vdd gnd cell_6t
Xbit_r53_c126 bl_126 br_126 wl_53 vdd gnd cell_6t
Xbit_r54_c126 bl_126 br_126 wl_54 vdd gnd cell_6t
Xbit_r55_c126 bl_126 br_126 wl_55 vdd gnd cell_6t
Xbit_r56_c126 bl_126 br_126 wl_56 vdd gnd cell_6t
Xbit_r57_c126 bl_126 br_126 wl_57 vdd gnd cell_6t
Xbit_r58_c126 bl_126 br_126 wl_58 vdd gnd cell_6t
Xbit_r59_c126 bl_126 br_126 wl_59 vdd gnd cell_6t
Xbit_r60_c126 bl_126 br_126 wl_60 vdd gnd cell_6t
Xbit_r61_c126 bl_126 br_126 wl_61 vdd gnd cell_6t
Xbit_r62_c126 bl_126 br_126 wl_62 vdd gnd cell_6t
Xbit_r63_c126 bl_126 br_126 wl_63 vdd gnd cell_6t
Xbit_r64_c126 bl_126 br_126 wl_64 vdd gnd cell_6t
Xbit_r65_c126 bl_126 br_126 wl_65 vdd gnd cell_6t
Xbit_r66_c126 bl_126 br_126 wl_66 vdd gnd cell_6t
Xbit_r67_c126 bl_126 br_126 wl_67 vdd gnd cell_6t
Xbit_r68_c126 bl_126 br_126 wl_68 vdd gnd cell_6t
Xbit_r69_c126 bl_126 br_126 wl_69 vdd gnd cell_6t
Xbit_r70_c126 bl_126 br_126 wl_70 vdd gnd cell_6t
Xbit_r71_c126 bl_126 br_126 wl_71 vdd gnd cell_6t
Xbit_r72_c126 bl_126 br_126 wl_72 vdd gnd cell_6t
Xbit_r73_c126 bl_126 br_126 wl_73 vdd gnd cell_6t
Xbit_r74_c126 bl_126 br_126 wl_74 vdd gnd cell_6t
Xbit_r75_c126 bl_126 br_126 wl_75 vdd gnd cell_6t
Xbit_r76_c126 bl_126 br_126 wl_76 vdd gnd cell_6t
Xbit_r77_c126 bl_126 br_126 wl_77 vdd gnd cell_6t
Xbit_r78_c126 bl_126 br_126 wl_78 vdd gnd cell_6t
Xbit_r79_c126 bl_126 br_126 wl_79 vdd gnd cell_6t
Xbit_r80_c126 bl_126 br_126 wl_80 vdd gnd cell_6t
Xbit_r81_c126 bl_126 br_126 wl_81 vdd gnd cell_6t
Xbit_r82_c126 bl_126 br_126 wl_82 vdd gnd cell_6t
Xbit_r83_c126 bl_126 br_126 wl_83 vdd gnd cell_6t
Xbit_r84_c126 bl_126 br_126 wl_84 vdd gnd cell_6t
Xbit_r85_c126 bl_126 br_126 wl_85 vdd gnd cell_6t
Xbit_r86_c126 bl_126 br_126 wl_86 vdd gnd cell_6t
Xbit_r87_c126 bl_126 br_126 wl_87 vdd gnd cell_6t
Xbit_r88_c126 bl_126 br_126 wl_88 vdd gnd cell_6t
Xbit_r89_c126 bl_126 br_126 wl_89 vdd gnd cell_6t
Xbit_r90_c126 bl_126 br_126 wl_90 vdd gnd cell_6t
Xbit_r91_c126 bl_126 br_126 wl_91 vdd gnd cell_6t
Xbit_r92_c126 bl_126 br_126 wl_92 vdd gnd cell_6t
Xbit_r93_c126 bl_126 br_126 wl_93 vdd gnd cell_6t
Xbit_r94_c126 bl_126 br_126 wl_94 vdd gnd cell_6t
Xbit_r95_c126 bl_126 br_126 wl_95 vdd gnd cell_6t
Xbit_r96_c126 bl_126 br_126 wl_96 vdd gnd cell_6t
Xbit_r97_c126 bl_126 br_126 wl_97 vdd gnd cell_6t
Xbit_r98_c126 bl_126 br_126 wl_98 vdd gnd cell_6t
Xbit_r99_c126 bl_126 br_126 wl_99 vdd gnd cell_6t
Xbit_r100_c126 bl_126 br_126 wl_100 vdd gnd cell_6t
Xbit_r101_c126 bl_126 br_126 wl_101 vdd gnd cell_6t
Xbit_r102_c126 bl_126 br_126 wl_102 vdd gnd cell_6t
Xbit_r103_c126 bl_126 br_126 wl_103 vdd gnd cell_6t
Xbit_r104_c126 bl_126 br_126 wl_104 vdd gnd cell_6t
Xbit_r105_c126 bl_126 br_126 wl_105 vdd gnd cell_6t
Xbit_r106_c126 bl_126 br_126 wl_106 vdd gnd cell_6t
Xbit_r107_c126 bl_126 br_126 wl_107 vdd gnd cell_6t
Xbit_r108_c126 bl_126 br_126 wl_108 vdd gnd cell_6t
Xbit_r109_c126 bl_126 br_126 wl_109 vdd gnd cell_6t
Xbit_r110_c126 bl_126 br_126 wl_110 vdd gnd cell_6t
Xbit_r111_c126 bl_126 br_126 wl_111 vdd gnd cell_6t
Xbit_r112_c126 bl_126 br_126 wl_112 vdd gnd cell_6t
Xbit_r113_c126 bl_126 br_126 wl_113 vdd gnd cell_6t
Xbit_r114_c126 bl_126 br_126 wl_114 vdd gnd cell_6t
Xbit_r115_c126 bl_126 br_126 wl_115 vdd gnd cell_6t
Xbit_r116_c126 bl_126 br_126 wl_116 vdd gnd cell_6t
Xbit_r117_c126 bl_126 br_126 wl_117 vdd gnd cell_6t
Xbit_r118_c126 bl_126 br_126 wl_118 vdd gnd cell_6t
Xbit_r119_c126 bl_126 br_126 wl_119 vdd gnd cell_6t
Xbit_r120_c126 bl_126 br_126 wl_120 vdd gnd cell_6t
Xbit_r121_c126 bl_126 br_126 wl_121 vdd gnd cell_6t
Xbit_r122_c126 bl_126 br_126 wl_122 vdd gnd cell_6t
Xbit_r123_c126 bl_126 br_126 wl_123 vdd gnd cell_6t
Xbit_r124_c126 bl_126 br_126 wl_124 vdd gnd cell_6t
Xbit_r125_c126 bl_126 br_126 wl_125 vdd gnd cell_6t
Xbit_r126_c126 bl_126 br_126 wl_126 vdd gnd cell_6t
Xbit_r127_c126 bl_126 br_126 wl_127 vdd gnd cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd cell_6t
Xbit_r1_c127 bl_127 br_127 wl_1 vdd gnd cell_6t
Xbit_r2_c127 bl_127 br_127 wl_2 vdd gnd cell_6t
Xbit_r3_c127 bl_127 br_127 wl_3 vdd gnd cell_6t
Xbit_r4_c127 bl_127 br_127 wl_4 vdd gnd cell_6t
Xbit_r5_c127 bl_127 br_127 wl_5 vdd gnd cell_6t
Xbit_r6_c127 bl_127 br_127 wl_6 vdd gnd cell_6t
Xbit_r7_c127 bl_127 br_127 wl_7 vdd gnd cell_6t
Xbit_r8_c127 bl_127 br_127 wl_8 vdd gnd cell_6t
Xbit_r9_c127 bl_127 br_127 wl_9 vdd gnd cell_6t
Xbit_r10_c127 bl_127 br_127 wl_10 vdd gnd cell_6t
Xbit_r11_c127 bl_127 br_127 wl_11 vdd gnd cell_6t
Xbit_r12_c127 bl_127 br_127 wl_12 vdd gnd cell_6t
Xbit_r13_c127 bl_127 br_127 wl_13 vdd gnd cell_6t
Xbit_r14_c127 bl_127 br_127 wl_14 vdd gnd cell_6t
Xbit_r15_c127 bl_127 br_127 wl_15 vdd gnd cell_6t
Xbit_r16_c127 bl_127 br_127 wl_16 vdd gnd cell_6t
Xbit_r17_c127 bl_127 br_127 wl_17 vdd gnd cell_6t
Xbit_r18_c127 bl_127 br_127 wl_18 vdd gnd cell_6t
Xbit_r19_c127 bl_127 br_127 wl_19 vdd gnd cell_6t
Xbit_r20_c127 bl_127 br_127 wl_20 vdd gnd cell_6t
Xbit_r21_c127 bl_127 br_127 wl_21 vdd gnd cell_6t
Xbit_r22_c127 bl_127 br_127 wl_22 vdd gnd cell_6t
Xbit_r23_c127 bl_127 br_127 wl_23 vdd gnd cell_6t
Xbit_r24_c127 bl_127 br_127 wl_24 vdd gnd cell_6t
Xbit_r25_c127 bl_127 br_127 wl_25 vdd gnd cell_6t
Xbit_r26_c127 bl_127 br_127 wl_26 vdd gnd cell_6t
Xbit_r27_c127 bl_127 br_127 wl_27 vdd gnd cell_6t
Xbit_r28_c127 bl_127 br_127 wl_28 vdd gnd cell_6t
Xbit_r29_c127 bl_127 br_127 wl_29 vdd gnd cell_6t
Xbit_r30_c127 bl_127 br_127 wl_30 vdd gnd cell_6t
Xbit_r31_c127 bl_127 br_127 wl_31 vdd gnd cell_6t
Xbit_r32_c127 bl_127 br_127 wl_32 vdd gnd cell_6t
Xbit_r33_c127 bl_127 br_127 wl_33 vdd gnd cell_6t
Xbit_r34_c127 bl_127 br_127 wl_34 vdd gnd cell_6t
Xbit_r35_c127 bl_127 br_127 wl_35 vdd gnd cell_6t
Xbit_r36_c127 bl_127 br_127 wl_36 vdd gnd cell_6t
Xbit_r37_c127 bl_127 br_127 wl_37 vdd gnd cell_6t
Xbit_r38_c127 bl_127 br_127 wl_38 vdd gnd cell_6t
Xbit_r39_c127 bl_127 br_127 wl_39 vdd gnd cell_6t
Xbit_r40_c127 bl_127 br_127 wl_40 vdd gnd cell_6t
Xbit_r41_c127 bl_127 br_127 wl_41 vdd gnd cell_6t
Xbit_r42_c127 bl_127 br_127 wl_42 vdd gnd cell_6t
Xbit_r43_c127 bl_127 br_127 wl_43 vdd gnd cell_6t
Xbit_r44_c127 bl_127 br_127 wl_44 vdd gnd cell_6t
Xbit_r45_c127 bl_127 br_127 wl_45 vdd gnd cell_6t
Xbit_r46_c127 bl_127 br_127 wl_46 vdd gnd cell_6t
Xbit_r47_c127 bl_127 br_127 wl_47 vdd gnd cell_6t
Xbit_r48_c127 bl_127 br_127 wl_48 vdd gnd cell_6t
Xbit_r49_c127 bl_127 br_127 wl_49 vdd gnd cell_6t
Xbit_r50_c127 bl_127 br_127 wl_50 vdd gnd cell_6t
Xbit_r51_c127 bl_127 br_127 wl_51 vdd gnd cell_6t
Xbit_r52_c127 bl_127 br_127 wl_52 vdd gnd cell_6t
Xbit_r53_c127 bl_127 br_127 wl_53 vdd gnd cell_6t
Xbit_r54_c127 bl_127 br_127 wl_54 vdd gnd cell_6t
Xbit_r55_c127 bl_127 br_127 wl_55 vdd gnd cell_6t
Xbit_r56_c127 bl_127 br_127 wl_56 vdd gnd cell_6t
Xbit_r57_c127 bl_127 br_127 wl_57 vdd gnd cell_6t
Xbit_r58_c127 bl_127 br_127 wl_58 vdd gnd cell_6t
Xbit_r59_c127 bl_127 br_127 wl_59 vdd gnd cell_6t
Xbit_r60_c127 bl_127 br_127 wl_60 vdd gnd cell_6t
Xbit_r61_c127 bl_127 br_127 wl_61 vdd gnd cell_6t
Xbit_r62_c127 bl_127 br_127 wl_62 vdd gnd cell_6t
Xbit_r63_c127 bl_127 br_127 wl_63 vdd gnd cell_6t
Xbit_r64_c127 bl_127 br_127 wl_64 vdd gnd cell_6t
Xbit_r65_c127 bl_127 br_127 wl_65 vdd gnd cell_6t
Xbit_r66_c127 bl_127 br_127 wl_66 vdd gnd cell_6t
Xbit_r67_c127 bl_127 br_127 wl_67 vdd gnd cell_6t
Xbit_r68_c127 bl_127 br_127 wl_68 vdd gnd cell_6t
Xbit_r69_c127 bl_127 br_127 wl_69 vdd gnd cell_6t
Xbit_r70_c127 bl_127 br_127 wl_70 vdd gnd cell_6t
Xbit_r71_c127 bl_127 br_127 wl_71 vdd gnd cell_6t
Xbit_r72_c127 bl_127 br_127 wl_72 vdd gnd cell_6t
Xbit_r73_c127 bl_127 br_127 wl_73 vdd gnd cell_6t
Xbit_r74_c127 bl_127 br_127 wl_74 vdd gnd cell_6t
Xbit_r75_c127 bl_127 br_127 wl_75 vdd gnd cell_6t
Xbit_r76_c127 bl_127 br_127 wl_76 vdd gnd cell_6t
Xbit_r77_c127 bl_127 br_127 wl_77 vdd gnd cell_6t
Xbit_r78_c127 bl_127 br_127 wl_78 vdd gnd cell_6t
Xbit_r79_c127 bl_127 br_127 wl_79 vdd gnd cell_6t
Xbit_r80_c127 bl_127 br_127 wl_80 vdd gnd cell_6t
Xbit_r81_c127 bl_127 br_127 wl_81 vdd gnd cell_6t
Xbit_r82_c127 bl_127 br_127 wl_82 vdd gnd cell_6t
Xbit_r83_c127 bl_127 br_127 wl_83 vdd gnd cell_6t
Xbit_r84_c127 bl_127 br_127 wl_84 vdd gnd cell_6t
Xbit_r85_c127 bl_127 br_127 wl_85 vdd gnd cell_6t
Xbit_r86_c127 bl_127 br_127 wl_86 vdd gnd cell_6t
Xbit_r87_c127 bl_127 br_127 wl_87 vdd gnd cell_6t
Xbit_r88_c127 bl_127 br_127 wl_88 vdd gnd cell_6t
Xbit_r89_c127 bl_127 br_127 wl_89 vdd gnd cell_6t
Xbit_r90_c127 bl_127 br_127 wl_90 vdd gnd cell_6t
Xbit_r91_c127 bl_127 br_127 wl_91 vdd gnd cell_6t
Xbit_r92_c127 bl_127 br_127 wl_92 vdd gnd cell_6t
Xbit_r93_c127 bl_127 br_127 wl_93 vdd gnd cell_6t
Xbit_r94_c127 bl_127 br_127 wl_94 vdd gnd cell_6t
Xbit_r95_c127 bl_127 br_127 wl_95 vdd gnd cell_6t
Xbit_r96_c127 bl_127 br_127 wl_96 vdd gnd cell_6t
Xbit_r97_c127 bl_127 br_127 wl_97 vdd gnd cell_6t
Xbit_r98_c127 bl_127 br_127 wl_98 vdd gnd cell_6t
Xbit_r99_c127 bl_127 br_127 wl_99 vdd gnd cell_6t
Xbit_r100_c127 bl_127 br_127 wl_100 vdd gnd cell_6t
Xbit_r101_c127 bl_127 br_127 wl_101 vdd gnd cell_6t
Xbit_r102_c127 bl_127 br_127 wl_102 vdd gnd cell_6t
Xbit_r103_c127 bl_127 br_127 wl_103 vdd gnd cell_6t
Xbit_r104_c127 bl_127 br_127 wl_104 vdd gnd cell_6t
Xbit_r105_c127 bl_127 br_127 wl_105 vdd gnd cell_6t
Xbit_r106_c127 bl_127 br_127 wl_106 vdd gnd cell_6t
Xbit_r107_c127 bl_127 br_127 wl_107 vdd gnd cell_6t
Xbit_r108_c127 bl_127 br_127 wl_108 vdd gnd cell_6t
Xbit_r109_c127 bl_127 br_127 wl_109 vdd gnd cell_6t
Xbit_r110_c127 bl_127 br_127 wl_110 vdd gnd cell_6t
Xbit_r111_c127 bl_127 br_127 wl_111 vdd gnd cell_6t
Xbit_r112_c127 bl_127 br_127 wl_112 vdd gnd cell_6t
Xbit_r113_c127 bl_127 br_127 wl_113 vdd gnd cell_6t
Xbit_r114_c127 bl_127 br_127 wl_114 vdd gnd cell_6t
Xbit_r115_c127 bl_127 br_127 wl_115 vdd gnd cell_6t
Xbit_r116_c127 bl_127 br_127 wl_116 vdd gnd cell_6t
Xbit_r117_c127 bl_127 br_127 wl_117 vdd gnd cell_6t
Xbit_r118_c127 bl_127 br_127 wl_118 vdd gnd cell_6t
Xbit_r119_c127 bl_127 br_127 wl_119 vdd gnd cell_6t
Xbit_r120_c127 bl_127 br_127 wl_120 vdd gnd cell_6t
Xbit_r121_c127 bl_127 br_127 wl_121 vdd gnd cell_6t
Xbit_r122_c127 bl_127 br_127 wl_122 vdd gnd cell_6t
Xbit_r123_c127 bl_127 br_127 wl_123 vdd gnd cell_6t
Xbit_r124_c127 bl_127 br_127 wl_124 vdd gnd cell_6t
Xbit_r125_c127 bl_127 br_127 wl_125 vdd gnd cell_6t
Xbit_r126_c127 bl_127 br_127 wl_126 vdd gnd cell_6t
Xbit_r127_c127 bl_127 br_127 wl_127 vdd gnd cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd cell_6t
Xbit_r1_c128 bl_128 br_128 wl_1 vdd gnd cell_6t
Xbit_r2_c128 bl_128 br_128 wl_2 vdd gnd cell_6t
Xbit_r3_c128 bl_128 br_128 wl_3 vdd gnd cell_6t
Xbit_r4_c128 bl_128 br_128 wl_4 vdd gnd cell_6t
Xbit_r5_c128 bl_128 br_128 wl_5 vdd gnd cell_6t
Xbit_r6_c128 bl_128 br_128 wl_6 vdd gnd cell_6t
Xbit_r7_c128 bl_128 br_128 wl_7 vdd gnd cell_6t
Xbit_r8_c128 bl_128 br_128 wl_8 vdd gnd cell_6t
Xbit_r9_c128 bl_128 br_128 wl_9 vdd gnd cell_6t
Xbit_r10_c128 bl_128 br_128 wl_10 vdd gnd cell_6t
Xbit_r11_c128 bl_128 br_128 wl_11 vdd gnd cell_6t
Xbit_r12_c128 bl_128 br_128 wl_12 vdd gnd cell_6t
Xbit_r13_c128 bl_128 br_128 wl_13 vdd gnd cell_6t
Xbit_r14_c128 bl_128 br_128 wl_14 vdd gnd cell_6t
Xbit_r15_c128 bl_128 br_128 wl_15 vdd gnd cell_6t
Xbit_r16_c128 bl_128 br_128 wl_16 vdd gnd cell_6t
Xbit_r17_c128 bl_128 br_128 wl_17 vdd gnd cell_6t
Xbit_r18_c128 bl_128 br_128 wl_18 vdd gnd cell_6t
Xbit_r19_c128 bl_128 br_128 wl_19 vdd gnd cell_6t
Xbit_r20_c128 bl_128 br_128 wl_20 vdd gnd cell_6t
Xbit_r21_c128 bl_128 br_128 wl_21 vdd gnd cell_6t
Xbit_r22_c128 bl_128 br_128 wl_22 vdd gnd cell_6t
Xbit_r23_c128 bl_128 br_128 wl_23 vdd gnd cell_6t
Xbit_r24_c128 bl_128 br_128 wl_24 vdd gnd cell_6t
Xbit_r25_c128 bl_128 br_128 wl_25 vdd gnd cell_6t
Xbit_r26_c128 bl_128 br_128 wl_26 vdd gnd cell_6t
Xbit_r27_c128 bl_128 br_128 wl_27 vdd gnd cell_6t
Xbit_r28_c128 bl_128 br_128 wl_28 vdd gnd cell_6t
Xbit_r29_c128 bl_128 br_128 wl_29 vdd gnd cell_6t
Xbit_r30_c128 bl_128 br_128 wl_30 vdd gnd cell_6t
Xbit_r31_c128 bl_128 br_128 wl_31 vdd gnd cell_6t
Xbit_r32_c128 bl_128 br_128 wl_32 vdd gnd cell_6t
Xbit_r33_c128 bl_128 br_128 wl_33 vdd gnd cell_6t
Xbit_r34_c128 bl_128 br_128 wl_34 vdd gnd cell_6t
Xbit_r35_c128 bl_128 br_128 wl_35 vdd gnd cell_6t
Xbit_r36_c128 bl_128 br_128 wl_36 vdd gnd cell_6t
Xbit_r37_c128 bl_128 br_128 wl_37 vdd gnd cell_6t
Xbit_r38_c128 bl_128 br_128 wl_38 vdd gnd cell_6t
Xbit_r39_c128 bl_128 br_128 wl_39 vdd gnd cell_6t
Xbit_r40_c128 bl_128 br_128 wl_40 vdd gnd cell_6t
Xbit_r41_c128 bl_128 br_128 wl_41 vdd gnd cell_6t
Xbit_r42_c128 bl_128 br_128 wl_42 vdd gnd cell_6t
Xbit_r43_c128 bl_128 br_128 wl_43 vdd gnd cell_6t
Xbit_r44_c128 bl_128 br_128 wl_44 vdd gnd cell_6t
Xbit_r45_c128 bl_128 br_128 wl_45 vdd gnd cell_6t
Xbit_r46_c128 bl_128 br_128 wl_46 vdd gnd cell_6t
Xbit_r47_c128 bl_128 br_128 wl_47 vdd gnd cell_6t
Xbit_r48_c128 bl_128 br_128 wl_48 vdd gnd cell_6t
Xbit_r49_c128 bl_128 br_128 wl_49 vdd gnd cell_6t
Xbit_r50_c128 bl_128 br_128 wl_50 vdd gnd cell_6t
Xbit_r51_c128 bl_128 br_128 wl_51 vdd gnd cell_6t
Xbit_r52_c128 bl_128 br_128 wl_52 vdd gnd cell_6t
Xbit_r53_c128 bl_128 br_128 wl_53 vdd gnd cell_6t
Xbit_r54_c128 bl_128 br_128 wl_54 vdd gnd cell_6t
Xbit_r55_c128 bl_128 br_128 wl_55 vdd gnd cell_6t
Xbit_r56_c128 bl_128 br_128 wl_56 vdd gnd cell_6t
Xbit_r57_c128 bl_128 br_128 wl_57 vdd gnd cell_6t
Xbit_r58_c128 bl_128 br_128 wl_58 vdd gnd cell_6t
Xbit_r59_c128 bl_128 br_128 wl_59 vdd gnd cell_6t
Xbit_r60_c128 bl_128 br_128 wl_60 vdd gnd cell_6t
Xbit_r61_c128 bl_128 br_128 wl_61 vdd gnd cell_6t
Xbit_r62_c128 bl_128 br_128 wl_62 vdd gnd cell_6t
Xbit_r63_c128 bl_128 br_128 wl_63 vdd gnd cell_6t
Xbit_r64_c128 bl_128 br_128 wl_64 vdd gnd cell_6t
Xbit_r65_c128 bl_128 br_128 wl_65 vdd gnd cell_6t
Xbit_r66_c128 bl_128 br_128 wl_66 vdd gnd cell_6t
Xbit_r67_c128 bl_128 br_128 wl_67 vdd gnd cell_6t
Xbit_r68_c128 bl_128 br_128 wl_68 vdd gnd cell_6t
Xbit_r69_c128 bl_128 br_128 wl_69 vdd gnd cell_6t
Xbit_r70_c128 bl_128 br_128 wl_70 vdd gnd cell_6t
Xbit_r71_c128 bl_128 br_128 wl_71 vdd gnd cell_6t
Xbit_r72_c128 bl_128 br_128 wl_72 vdd gnd cell_6t
Xbit_r73_c128 bl_128 br_128 wl_73 vdd gnd cell_6t
Xbit_r74_c128 bl_128 br_128 wl_74 vdd gnd cell_6t
Xbit_r75_c128 bl_128 br_128 wl_75 vdd gnd cell_6t
Xbit_r76_c128 bl_128 br_128 wl_76 vdd gnd cell_6t
Xbit_r77_c128 bl_128 br_128 wl_77 vdd gnd cell_6t
Xbit_r78_c128 bl_128 br_128 wl_78 vdd gnd cell_6t
Xbit_r79_c128 bl_128 br_128 wl_79 vdd gnd cell_6t
Xbit_r80_c128 bl_128 br_128 wl_80 vdd gnd cell_6t
Xbit_r81_c128 bl_128 br_128 wl_81 vdd gnd cell_6t
Xbit_r82_c128 bl_128 br_128 wl_82 vdd gnd cell_6t
Xbit_r83_c128 bl_128 br_128 wl_83 vdd gnd cell_6t
Xbit_r84_c128 bl_128 br_128 wl_84 vdd gnd cell_6t
Xbit_r85_c128 bl_128 br_128 wl_85 vdd gnd cell_6t
Xbit_r86_c128 bl_128 br_128 wl_86 vdd gnd cell_6t
Xbit_r87_c128 bl_128 br_128 wl_87 vdd gnd cell_6t
Xbit_r88_c128 bl_128 br_128 wl_88 vdd gnd cell_6t
Xbit_r89_c128 bl_128 br_128 wl_89 vdd gnd cell_6t
Xbit_r90_c128 bl_128 br_128 wl_90 vdd gnd cell_6t
Xbit_r91_c128 bl_128 br_128 wl_91 vdd gnd cell_6t
Xbit_r92_c128 bl_128 br_128 wl_92 vdd gnd cell_6t
Xbit_r93_c128 bl_128 br_128 wl_93 vdd gnd cell_6t
Xbit_r94_c128 bl_128 br_128 wl_94 vdd gnd cell_6t
Xbit_r95_c128 bl_128 br_128 wl_95 vdd gnd cell_6t
Xbit_r96_c128 bl_128 br_128 wl_96 vdd gnd cell_6t
Xbit_r97_c128 bl_128 br_128 wl_97 vdd gnd cell_6t
Xbit_r98_c128 bl_128 br_128 wl_98 vdd gnd cell_6t
Xbit_r99_c128 bl_128 br_128 wl_99 vdd gnd cell_6t
Xbit_r100_c128 bl_128 br_128 wl_100 vdd gnd cell_6t
Xbit_r101_c128 bl_128 br_128 wl_101 vdd gnd cell_6t
Xbit_r102_c128 bl_128 br_128 wl_102 vdd gnd cell_6t
Xbit_r103_c128 bl_128 br_128 wl_103 vdd gnd cell_6t
Xbit_r104_c128 bl_128 br_128 wl_104 vdd gnd cell_6t
Xbit_r105_c128 bl_128 br_128 wl_105 vdd gnd cell_6t
Xbit_r106_c128 bl_128 br_128 wl_106 vdd gnd cell_6t
Xbit_r107_c128 bl_128 br_128 wl_107 vdd gnd cell_6t
Xbit_r108_c128 bl_128 br_128 wl_108 vdd gnd cell_6t
Xbit_r109_c128 bl_128 br_128 wl_109 vdd gnd cell_6t
Xbit_r110_c128 bl_128 br_128 wl_110 vdd gnd cell_6t
Xbit_r111_c128 bl_128 br_128 wl_111 vdd gnd cell_6t
Xbit_r112_c128 bl_128 br_128 wl_112 vdd gnd cell_6t
Xbit_r113_c128 bl_128 br_128 wl_113 vdd gnd cell_6t
Xbit_r114_c128 bl_128 br_128 wl_114 vdd gnd cell_6t
Xbit_r115_c128 bl_128 br_128 wl_115 vdd gnd cell_6t
Xbit_r116_c128 bl_128 br_128 wl_116 vdd gnd cell_6t
Xbit_r117_c128 bl_128 br_128 wl_117 vdd gnd cell_6t
Xbit_r118_c128 bl_128 br_128 wl_118 vdd gnd cell_6t
Xbit_r119_c128 bl_128 br_128 wl_119 vdd gnd cell_6t
Xbit_r120_c128 bl_128 br_128 wl_120 vdd gnd cell_6t
Xbit_r121_c128 bl_128 br_128 wl_121 vdd gnd cell_6t
Xbit_r122_c128 bl_128 br_128 wl_122 vdd gnd cell_6t
Xbit_r123_c128 bl_128 br_128 wl_123 vdd gnd cell_6t
Xbit_r124_c128 bl_128 br_128 wl_124 vdd gnd cell_6t
Xbit_r125_c128 bl_128 br_128 wl_125 vdd gnd cell_6t
Xbit_r126_c128 bl_128 br_128 wl_126 vdd gnd cell_6t
Xbit_r127_c128 bl_128 br_128 wl_127 vdd gnd cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd cell_6t
Xbit_r1_c129 bl_129 br_129 wl_1 vdd gnd cell_6t
Xbit_r2_c129 bl_129 br_129 wl_2 vdd gnd cell_6t
Xbit_r3_c129 bl_129 br_129 wl_3 vdd gnd cell_6t
Xbit_r4_c129 bl_129 br_129 wl_4 vdd gnd cell_6t
Xbit_r5_c129 bl_129 br_129 wl_5 vdd gnd cell_6t
Xbit_r6_c129 bl_129 br_129 wl_6 vdd gnd cell_6t
Xbit_r7_c129 bl_129 br_129 wl_7 vdd gnd cell_6t
Xbit_r8_c129 bl_129 br_129 wl_8 vdd gnd cell_6t
Xbit_r9_c129 bl_129 br_129 wl_9 vdd gnd cell_6t
Xbit_r10_c129 bl_129 br_129 wl_10 vdd gnd cell_6t
Xbit_r11_c129 bl_129 br_129 wl_11 vdd gnd cell_6t
Xbit_r12_c129 bl_129 br_129 wl_12 vdd gnd cell_6t
Xbit_r13_c129 bl_129 br_129 wl_13 vdd gnd cell_6t
Xbit_r14_c129 bl_129 br_129 wl_14 vdd gnd cell_6t
Xbit_r15_c129 bl_129 br_129 wl_15 vdd gnd cell_6t
Xbit_r16_c129 bl_129 br_129 wl_16 vdd gnd cell_6t
Xbit_r17_c129 bl_129 br_129 wl_17 vdd gnd cell_6t
Xbit_r18_c129 bl_129 br_129 wl_18 vdd gnd cell_6t
Xbit_r19_c129 bl_129 br_129 wl_19 vdd gnd cell_6t
Xbit_r20_c129 bl_129 br_129 wl_20 vdd gnd cell_6t
Xbit_r21_c129 bl_129 br_129 wl_21 vdd gnd cell_6t
Xbit_r22_c129 bl_129 br_129 wl_22 vdd gnd cell_6t
Xbit_r23_c129 bl_129 br_129 wl_23 vdd gnd cell_6t
Xbit_r24_c129 bl_129 br_129 wl_24 vdd gnd cell_6t
Xbit_r25_c129 bl_129 br_129 wl_25 vdd gnd cell_6t
Xbit_r26_c129 bl_129 br_129 wl_26 vdd gnd cell_6t
Xbit_r27_c129 bl_129 br_129 wl_27 vdd gnd cell_6t
Xbit_r28_c129 bl_129 br_129 wl_28 vdd gnd cell_6t
Xbit_r29_c129 bl_129 br_129 wl_29 vdd gnd cell_6t
Xbit_r30_c129 bl_129 br_129 wl_30 vdd gnd cell_6t
Xbit_r31_c129 bl_129 br_129 wl_31 vdd gnd cell_6t
Xbit_r32_c129 bl_129 br_129 wl_32 vdd gnd cell_6t
Xbit_r33_c129 bl_129 br_129 wl_33 vdd gnd cell_6t
Xbit_r34_c129 bl_129 br_129 wl_34 vdd gnd cell_6t
Xbit_r35_c129 bl_129 br_129 wl_35 vdd gnd cell_6t
Xbit_r36_c129 bl_129 br_129 wl_36 vdd gnd cell_6t
Xbit_r37_c129 bl_129 br_129 wl_37 vdd gnd cell_6t
Xbit_r38_c129 bl_129 br_129 wl_38 vdd gnd cell_6t
Xbit_r39_c129 bl_129 br_129 wl_39 vdd gnd cell_6t
Xbit_r40_c129 bl_129 br_129 wl_40 vdd gnd cell_6t
Xbit_r41_c129 bl_129 br_129 wl_41 vdd gnd cell_6t
Xbit_r42_c129 bl_129 br_129 wl_42 vdd gnd cell_6t
Xbit_r43_c129 bl_129 br_129 wl_43 vdd gnd cell_6t
Xbit_r44_c129 bl_129 br_129 wl_44 vdd gnd cell_6t
Xbit_r45_c129 bl_129 br_129 wl_45 vdd gnd cell_6t
Xbit_r46_c129 bl_129 br_129 wl_46 vdd gnd cell_6t
Xbit_r47_c129 bl_129 br_129 wl_47 vdd gnd cell_6t
Xbit_r48_c129 bl_129 br_129 wl_48 vdd gnd cell_6t
Xbit_r49_c129 bl_129 br_129 wl_49 vdd gnd cell_6t
Xbit_r50_c129 bl_129 br_129 wl_50 vdd gnd cell_6t
Xbit_r51_c129 bl_129 br_129 wl_51 vdd gnd cell_6t
Xbit_r52_c129 bl_129 br_129 wl_52 vdd gnd cell_6t
Xbit_r53_c129 bl_129 br_129 wl_53 vdd gnd cell_6t
Xbit_r54_c129 bl_129 br_129 wl_54 vdd gnd cell_6t
Xbit_r55_c129 bl_129 br_129 wl_55 vdd gnd cell_6t
Xbit_r56_c129 bl_129 br_129 wl_56 vdd gnd cell_6t
Xbit_r57_c129 bl_129 br_129 wl_57 vdd gnd cell_6t
Xbit_r58_c129 bl_129 br_129 wl_58 vdd gnd cell_6t
Xbit_r59_c129 bl_129 br_129 wl_59 vdd gnd cell_6t
Xbit_r60_c129 bl_129 br_129 wl_60 vdd gnd cell_6t
Xbit_r61_c129 bl_129 br_129 wl_61 vdd gnd cell_6t
Xbit_r62_c129 bl_129 br_129 wl_62 vdd gnd cell_6t
Xbit_r63_c129 bl_129 br_129 wl_63 vdd gnd cell_6t
Xbit_r64_c129 bl_129 br_129 wl_64 vdd gnd cell_6t
Xbit_r65_c129 bl_129 br_129 wl_65 vdd gnd cell_6t
Xbit_r66_c129 bl_129 br_129 wl_66 vdd gnd cell_6t
Xbit_r67_c129 bl_129 br_129 wl_67 vdd gnd cell_6t
Xbit_r68_c129 bl_129 br_129 wl_68 vdd gnd cell_6t
Xbit_r69_c129 bl_129 br_129 wl_69 vdd gnd cell_6t
Xbit_r70_c129 bl_129 br_129 wl_70 vdd gnd cell_6t
Xbit_r71_c129 bl_129 br_129 wl_71 vdd gnd cell_6t
Xbit_r72_c129 bl_129 br_129 wl_72 vdd gnd cell_6t
Xbit_r73_c129 bl_129 br_129 wl_73 vdd gnd cell_6t
Xbit_r74_c129 bl_129 br_129 wl_74 vdd gnd cell_6t
Xbit_r75_c129 bl_129 br_129 wl_75 vdd gnd cell_6t
Xbit_r76_c129 bl_129 br_129 wl_76 vdd gnd cell_6t
Xbit_r77_c129 bl_129 br_129 wl_77 vdd gnd cell_6t
Xbit_r78_c129 bl_129 br_129 wl_78 vdd gnd cell_6t
Xbit_r79_c129 bl_129 br_129 wl_79 vdd gnd cell_6t
Xbit_r80_c129 bl_129 br_129 wl_80 vdd gnd cell_6t
Xbit_r81_c129 bl_129 br_129 wl_81 vdd gnd cell_6t
Xbit_r82_c129 bl_129 br_129 wl_82 vdd gnd cell_6t
Xbit_r83_c129 bl_129 br_129 wl_83 vdd gnd cell_6t
Xbit_r84_c129 bl_129 br_129 wl_84 vdd gnd cell_6t
Xbit_r85_c129 bl_129 br_129 wl_85 vdd gnd cell_6t
Xbit_r86_c129 bl_129 br_129 wl_86 vdd gnd cell_6t
Xbit_r87_c129 bl_129 br_129 wl_87 vdd gnd cell_6t
Xbit_r88_c129 bl_129 br_129 wl_88 vdd gnd cell_6t
Xbit_r89_c129 bl_129 br_129 wl_89 vdd gnd cell_6t
Xbit_r90_c129 bl_129 br_129 wl_90 vdd gnd cell_6t
Xbit_r91_c129 bl_129 br_129 wl_91 vdd gnd cell_6t
Xbit_r92_c129 bl_129 br_129 wl_92 vdd gnd cell_6t
Xbit_r93_c129 bl_129 br_129 wl_93 vdd gnd cell_6t
Xbit_r94_c129 bl_129 br_129 wl_94 vdd gnd cell_6t
Xbit_r95_c129 bl_129 br_129 wl_95 vdd gnd cell_6t
Xbit_r96_c129 bl_129 br_129 wl_96 vdd gnd cell_6t
Xbit_r97_c129 bl_129 br_129 wl_97 vdd gnd cell_6t
Xbit_r98_c129 bl_129 br_129 wl_98 vdd gnd cell_6t
Xbit_r99_c129 bl_129 br_129 wl_99 vdd gnd cell_6t
Xbit_r100_c129 bl_129 br_129 wl_100 vdd gnd cell_6t
Xbit_r101_c129 bl_129 br_129 wl_101 vdd gnd cell_6t
Xbit_r102_c129 bl_129 br_129 wl_102 vdd gnd cell_6t
Xbit_r103_c129 bl_129 br_129 wl_103 vdd gnd cell_6t
Xbit_r104_c129 bl_129 br_129 wl_104 vdd gnd cell_6t
Xbit_r105_c129 bl_129 br_129 wl_105 vdd gnd cell_6t
Xbit_r106_c129 bl_129 br_129 wl_106 vdd gnd cell_6t
Xbit_r107_c129 bl_129 br_129 wl_107 vdd gnd cell_6t
Xbit_r108_c129 bl_129 br_129 wl_108 vdd gnd cell_6t
Xbit_r109_c129 bl_129 br_129 wl_109 vdd gnd cell_6t
Xbit_r110_c129 bl_129 br_129 wl_110 vdd gnd cell_6t
Xbit_r111_c129 bl_129 br_129 wl_111 vdd gnd cell_6t
Xbit_r112_c129 bl_129 br_129 wl_112 vdd gnd cell_6t
Xbit_r113_c129 bl_129 br_129 wl_113 vdd gnd cell_6t
Xbit_r114_c129 bl_129 br_129 wl_114 vdd gnd cell_6t
Xbit_r115_c129 bl_129 br_129 wl_115 vdd gnd cell_6t
Xbit_r116_c129 bl_129 br_129 wl_116 vdd gnd cell_6t
Xbit_r117_c129 bl_129 br_129 wl_117 vdd gnd cell_6t
Xbit_r118_c129 bl_129 br_129 wl_118 vdd gnd cell_6t
Xbit_r119_c129 bl_129 br_129 wl_119 vdd gnd cell_6t
Xbit_r120_c129 bl_129 br_129 wl_120 vdd gnd cell_6t
Xbit_r121_c129 bl_129 br_129 wl_121 vdd gnd cell_6t
Xbit_r122_c129 bl_129 br_129 wl_122 vdd gnd cell_6t
Xbit_r123_c129 bl_129 br_129 wl_123 vdd gnd cell_6t
Xbit_r124_c129 bl_129 br_129 wl_124 vdd gnd cell_6t
Xbit_r125_c129 bl_129 br_129 wl_125 vdd gnd cell_6t
Xbit_r126_c129 bl_129 br_129 wl_126 vdd gnd cell_6t
Xbit_r127_c129 bl_129 br_129 wl_127 vdd gnd cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd cell_6t
Xbit_r1_c130 bl_130 br_130 wl_1 vdd gnd cell_6t
Xbit_r2_c130 bl_130 br_130 wl_2 vdd gnd cell_6t
Xbit_r3_c130 bl_130 br_130 wl_3 vdd gnd cell_6t
Xbit_r4_c130 bl_130 br_130 wl_4 vdd gnd cell_6t
Xbit_r5_c130 bl_130 br_130 wl_5 vdd gnd cell_6t
Xbit_r6_c130 bl_130 br_130 wl_6 vdd gnd cell_6t
Xbit_r7_c130 bl_130 br_130 wl_7 vdd gnd cell_6t
Xbit_r8_c130 bl_130 br_130 wl_8 vdd gnd cell_6t
Xbit_r9_c130 bl_130 br_130 wl_9 vdd gnd cell_6t
Xbit_r10_c130 bl_130 br_130 wl_10 vdd gnd cell_6t
Xbit_r11_c130 bl_130 br_130 wl_11 vdd gnd cell_6t
Xbit_r12_c130 bl_130 br_130 wl_12 vdd gnd cell_6t
Xbit_r13_c130 bl_130 br_130 wl_13 vdd gnd cell_6t
Xbit_r14_c130 bl_130 br_130 wl_14 vdd gnd cell_6t
Xbit_r15_c130 bl_130 br_130 wl_15 vdd gnd cell_6t
Xbit_r16_c130 bl_130 br_130 wl_16 vdd gnd cell_6t
Xbit_r17_c130 bl_130 br_130 wl_17 vdd gnd cell_6t
Xbit_r18_c130 bl_130 br_130 wl_18 vdd gnd cell_6t
Xbit_r19_c130 bl_130 br_130 wl_19 vdd gnd cell_6t
Xbit_r20_c130 bl_130 br_130 wl_20 vdd gnd cell_6t
Xbit_r21_c130 bl_130 br_130 wl_21 vdd gnd cell_6t
Xbit_r22_c130 bl_130 br_130 wl_22 vdd gnd cell_6t
Xbit_r23_c130 bl_130 br_130 wl_23 vdd gnd cell_6t
Xbit_r24_c130 bl_130 br_130 wl_24 vdd gnd cell_6t
Xbit_r25_c130 bl_130 br_130 wl_25 vdd gnd cell_6t
Xbit_r26_c130 bl_130 br_130 wl_26 vdd gnd cell_6t
Xbit_r27_c130 bl_130 br_130 wl_27 vdd gnd cell_6t
Xbit_r28_c130 bl_130 br_130 wl_28 vdd gnd cell_6t
Xbit_r29_c130 bl_130 br_130 wl_29 vdd gnd cell_6t
Xbit_r30_c130 bl_130 br_130 wl_30 vdd gnd cell_6t
Xbit_r31_c130 bl_130 br_130 wl_31 vdd gnd cell_6t
Xbit_r32_c130 bl_130 br_130 wl_32 vdd gnd cell_6t
Xbit_r33_c130 bl_130 br_130 wl_33 vdd gnd cell_6t
Xbit_r34_c130 bl_130 br_130 wl_34 vdd gnd cell_6t
Xbit_r35_c130 bl_130 br_130 wl_35 vdd gnd cell_6t
Xbit_r36_c130 bl_130 br_130 wl_36 vdd gnd cell_6t
Xbit_r37_c130 bl_130 br_130 wl_37 vdd gnd cell_6t
Xbit_r38_c130 bl_130 br_130 wl_38 vdd gnd cell_6t
Xbit_r39_c130 bl_130 br_130 wl_39 vdd gnd cell_6t
Xbit_r40_c130 bl_130 br_130 wl_40 vdd gnd cell_6t
Xbit_r41_c130 bl_130 br_130 wl_41 vdd gnd cell_6t
Xbit_r42_c130 bl_130 br_130 wl_42 vdd gnd cell_6t
Xbit_r43_c130 bl_130 br_130 wl_43 vdd gnd cell_6t
Xbit_r44_c130 bl_130 br_130 wl_44 vdd gnd cell_6t
Xbit_r45_c130 bl_130 br_130 wl_45 vdd gnd cell_6t
Xbit_r46_c130 bl_130 br_130 wl_46 vdd gnd cell_6t
Xbit_r47_c130 bl_130 br_130 wl_47 vdd gnd cell_6t
Xbit_r48_c130 bl_130 br_130 wl_48 vdd gnd cell_6t
Xbit_r49_c130 bl_130 br_130 wl_49 vdd gnd cell_6t
Xbit_r50_c130 bl_130 br_130 wl_50 vdd gnd cell_6t
Xbit_r51_c130 bl_130 br_130 wl_51 vdd gnd cell_6t
Xbit_r52_c130 bl_130 br_130 wl_52 vdd gnd cell_6t
Xbit_r53_c130 bl_130 br_130 wl_53 vdd gnd cell_6t
Xbit_r54_c130 bl_130 br_130 wl_54 vdd gnd cell_6t
Xbit_r55_c130 bl_130 br_130 wl_55 vdd gnd cell_6t
Xbit_r56_c130 bl_130 br_130 wl_56 vdd gnd cell_6t
Xbit_r57_c130 bl_130 br_130 wl_57 vdd gnd cell_6t
Xbit_r58_c130 bl_130 br_130 wl_58 vdd gnd cell_6t
Xbit_r59_c130 bl_130 br_130 wl_59 vdd gnd cell_6t
Xbit_r60_c130 bl_130 br_130 wl_60 vdd gnd cell_6t
Xbit_r61_c130 bl_130 br_130 wl_61 vdd gnd cell_6t
Xbit_r62_c130 bl_130 br_130 wl_62 vdd gnd cell_6t
Xbit_r63_c130 bl_130 br_130 wl_63 vdd gnd cell_6t
Xbit_r64_c130 bl_130 br_130 wl_64 vdd gnd cell_6t
Xbit_r65_c130 bl_130 br_130 wl_65 vdd gnd cell_6t
Xbit_r66_c130 bl_130 br_130 wl_66 vdd gnd cell_6t
Xbit_r67_c130 bl_130 br_130 wl_67 vdd gnd cell_6t
Xbit_r68_c130 bl_130 br_130 wl_68 vdd gnd cell_6t
Xbit_r69_c130 bl_130 br_130 wl_69 vdd gnd cell_6t
Xbit_r70_c130 bl_130 br_130 wl_70 vdd gnd cell_6t
Xbit_r71_c130 bl_130 br_130 wl_71 vdd gnd cell_6t
Xbit_r72_c130 bl_130 br_130 wl_72 vdd gnd cell_6t
Xbit_r73_c130 bl_130 br_130 wl_73 vdd gnd cell_6t
Xbit_r74_c130 bl_130 br_130 wl_74 vdd gnd cell_6t
Xbit_r75_c130 bl_130 br_130 wl_75 vdd gnd cell_6t
Xbit_r76_c130 bl_130 br_130 wl_76 vdd gnd cell_6t
Xbit_r77_c130 bl_130 br_130 wl_77 vdd gnd cell_6t
Xbit_r78_c130 bl_130 br_130 wl_78 vdd gnd cell_6t
Xbit_r79_c130 bl_130 br_130 wl_79 vdd gnd cell_6t
Xbit_r80_c130 bl_130 br_130 wl_80 vdd gnd cell_6t
Xbit_r81_c130 bl_130 br_130 wl_81 vdd gnd cell_6t
Xbit_r82_c130 bl_130 br_130 wl_82 vdd gnd cell_6t
Xbit_r83_c130 bl_130 br_130 wl_83 vdd gnd cell_6t
Xbit_r84_c130 bl_130 br_130 wl_84 vdd gnd cell_6t
Xbit_r85_c130 bl_130 br_130 wl_85 vdd gnd cell_6t
Xbit_r86_c130 bl_130 br_130 wl_86 vdd gnd cell_6t
Xbit_r87_c130 bl_130 br_130 wl_87 vdd gnd cell_6t
Xbit_r88_c130 bl_130 br_130 wl_88 vdd gnd cell_6t
Xbit_r89_c130 bl_130 br_130 wl_89 vdd gnd cell_6t
Xbit_r90_c130 bl_130 br_130 wl_90 vdd gnd cell_6t
Xbit_r91_c130 bl_130 br_130 wl_91 vdd gnd cell_6t
Xbit_r92_c130 bl_130 br_130 wl_92 vdd gnd cell_6t
Xbit_r93_c130 bl_130 br_130 wl_93 vdd gnd cell_6t
Xbit_r94_c130 bl_130 br_130 wl_94 vdd gnd cell_6t
Xbit_r95_c130 bl_130 br_130 wl_95 vdd gnd cell_6t
Xbit_r96_c130 bl_130 br_130 wl_96 vdd gnd cell_6t
Xbit_r97_c130 bl_130 br_130 wl_97 vdd gnd cell_6t
Xbit_r98_c130 bl_130 br_130 wl_98 vdd gnd cell_6t
Xbit_r99_c130 bl_130 br_130 wl_99 vdd gnd cell_6t
Xbit_r100_c130 bl_130 br_130 wl_100 vdd gnd cell_6t
Xbit_r101_c130 bl_130 br_130 wl_101 vdd gnd cell_6t
Xbit_r102_c130 bl_130 br_130 wl_102 vdd gnd cell_6t
Xbit_r103_c130 bl_130 br_130 wl_103 vdd gnd cell_6t
Xbit_r104_c130 bl_130 br_130 wl_104 vdd gnd cell_6t
Xbit_r105_c130 bl_130 br_130 wl_105 vdd gnd cell_6t
Xbit_r106_c130 bl_130 br_130 wl_106 vdd gnd cell_6t
Xbit_r107_c130 bl_130 br_130 wl_107 vdd gnd cell_6t
Xbit_r108_c130 bl_130 br_130 wl_108 vdd gnd cell_6t
Xbit_r109_c130 bl_130 br_130 wl_109 vdd gnd cell_6t
Xbit_r110_c130 bl_130 br_130 wl_110 vdd gnd cell_6t
Xbit_r111_c130 bl_130 br_130 wl_111 vdd gnd cell_6t
Xbit_r112_c130 bl_130 br_130 wl_112 vdd gnd cell_6t
Xbit_r113_c130 bl_130 br_130 wl_113 vdd gnd cell_6t
Xbit_r114_c130 bl_130 br_130 wl_114 vdd gnd cell_6t
Xbit_r115_c130 bl_130 br_130 wl_115 vdd gnd cell_6t
Xbit_r116_c130 bl_130 br_130 wl_116 vdd gnd cell_6t
Xbit_r117_c130 bl_130 br_130 wl_117 vdd gnd cell_6t
Xbit_r118_c130 bl_130 br_130 wl_118 vdd gnd cell_6t
Xbit_r119_c130 bl_130 br_130 wl_119 vdd gnd cell_6t
Xbit_r120_c130 bl_130 br_130 wl_120 vdd gnd cell_6t
Xbit_r121_c130 bl_130 br_130 wl_121 vdd gnd cell_6t
Xbit_r122_c130 bl_130 br_130 wl_122 vdd gnd cell_6t
Xbit_r123_c130 bl_130 br_130 wl_123 vdd gnd cell_6t
Xbit_r124_c130 bl_130 br_130 wl_124 vdd gnd cell_6t
Xbit_r125_c130 bl_130 br_130 wl_125 vdd gnd cell_6t
Xbit_r126_c130 bl_130 br_130 wl_126 vdd gnd cell_6t
Xbit_r127_c130 bl_130 br_130 wl_127 vdd gnd cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd cell_6t
Xbit_r1_c131 bl_131 br_131 wl_1 vdd gnd cell_6t
Xbit_r2_c131 bl_131 br_131 wl_2 vdd gnd cell_6t
Xbit_r3_c131 bl_131 br_131 wl_3 vdd gnd cell_6t
Xbit_r4_c131 bl_131 br_131 wl_4 vdd gnd cell_6t
Xbit_r5_c131 bl_131 br_131 wl_5 vdd gnd cell_6t
Xbit_r6_c131 bl_131 br_131 wl_6 vdd gnd cell_6t
Xbit_r7_c131 bl_131 br_131 wl_7 vdd gnd cell_6t
Xbit_r8_c131 bl_131 br_131 wl_8 vdd gnd cell_6t
Xbit_r9_c131 bl_131 br_131 wl_9 vdd gnd cell_6t
Xbit_r10_c131 bl_131 br_131 wl_10 vdd gnd cell_6t
Xbit_r11_c131 bl_131 br_131 wl_11 vdd gnd cell_6t
Xbit_r12_c131 bl_131 br_131 wl_12 vdd gnd cell_6t
Xbit_r13_c131 bl_131 br_131 wl_13 vdd gnd cell_6t
Xbit_r14_c131 bl_131 br_131 wl_14 vdd gnd cell_6t
Xbit_r15_c131 bl_131 br_131 wl_15 vdd gnd cell_6t
Xbit_r16_c131 bl_131 br_131 wl_16 vdd gnd cell_6t
Xbit_r17_c131 bl_131 br_131 wl_17 vdd gnd cell_6t
Xbit_r18_c131 bl_131 br_131 wl_18 vdd gnd cell_6t
Xbit_r19_c131 bl_131 br_131 wl_19 vdd gnd cell_6t
Xbit_r20_c131 bl_131 br_131 wl_20 vdd gnd cell_6t
Xbit_r21_c131 bl_131 br_131 wl_21 vdd gnd cell_6t
Xbit_r22_c131 bl_131 br_131 wl_22 vdd gnd cell_6t
Xbit_r23_c131 bl_131 br_131 wl_23 vdd gnd cell_6t
Xbit_r24_c131 bl_131 br_131 wl_24 vdd gnd cell_6t
Xbit_r25_c131 bl_131 br_131 wl_25 vdd gnd cell_6t
Xbit_r26_c131 bl_131 br_131 wl_26 vdd gnd cell_6t
Xbit_r27_c131 bl_131 br_131 wl_27 vdd gnd cell_6t
Xbit_r28_c131 bl_131 br_131 wl_28 vdd gnd cell_6t
Xbit_r29_c131 bl_131 br_131 wl_29 vdd gnd cell_6t
Xbit_r30_c131 bl_131 br_131 wl_30 vdd gnd cell_6t
Xbit_r31_c131 bl_131 br_131 wl_31 vdd gnd cell_6t
Xbit_r32_c131 bl_131 br_131 wl_32 vdd gnd cell_6t
Xbit_r33_c131 bl_131 br_131 wl_33 vdd gnd cell_6t
Xbit_r34_c131 bl_131 br_131 wl_34 vdd gnd cell_6t
Xbit_r35_c131 bl_131 br_131 wl_35 vdd gnd cell_6t
Xbit_r36_c131 bl_131 br_131 wl_36 vdd gnd cell_6t
Xbit_r37_c131 bl_131 br_131 wl_37 vdd gnd cell_6t
Xbit_r38_c131 bl_131 br_131 wl_38 vdd gnd cell_6t
Xbit_r39_c131 bl_131 br_131 wl_39 vdd gnd cell_6t
Xbit_r40_c131 bl_131 br_131 wl_40 vdd gnd cell_6t
Xbit_r41_c131 bl_131 br_131 wl_41 vdd gnd cell_6t
Xbit_r42_c131 bl_131 br_131 wl_42 vdd gnd cell_6t
Xbit_r43_c131 bl_131 br_131 wl_43 vdd gnd cell_6t
Xbit_r44_c131 bl_131 br_131 wl_44 vdd gnd cell_6t
Xbit_r45_c131 bl_131 br_131 wl_45 vdd gnd cell_6t
Xbit_r46_c131 bl_131 br_131 wl_46 vdd gnd cell_6t
Xbit_r47_c131 bl_131 br_131 wl_47 vdd gnd cell_6t
Xbit_r48_c131 bl_131 br_131 wl_48 vdd gnd cell_6t
Xbit_r49_c131 bl_131 br_131 wl_49 vdd gnd cell_6t
Xbit_r50_c131 bl_131 br_131 wl_50 vdd gnd cell_6t
Xbit_r51_c131 bl_131 br_131 wl_51 vdd gnd cell_6t
Xbit_r52_c131 bl_131 br_131 wl_52 vdd gnd cell_6t
Xbit_r53_c131 bl_131 br_131 wl_53 vdd gnd cell_6t
Xbit_r54_c131 bl_131 br_131 wl_54 vdd gnd cell_6t
Xbit_r55_c131 bl_131 br_131 wl_55 vdd gnd cell_6t
Xbit_r56_c131 bl_131 br_131 wl_56 vdd gnd cell_6t
Xbit_r57_c131 bl_131 br_131 wl_57 vdd gnd cell_6t
Xbit_r58_c131 bl_131 br_131 wl_58 vdd gnd cell_6t
Xbit_r59_c131 bl_131 br_131 wl_59 vdd gnd cell_6t
Xbit_r60_c131 bl_131 br_131 wl_60 vdd gnd cell_6t
Xbit_r61_c131 bl_131 br_131 wl_61 vdd gnd cell_6t
Xbit_r62_c131 bl_131 br_131 wl_62 vdd gnd cell_6t
Xbit_r63_c131 bl_131 br_131 wl_63 vdd gnd cell_6t
Xbit_r64_c131 bl_131 br_131 wl_64 vdd gnd cell_6t
Xbit_r65_c131 bl_131 br_131 wl_65 vdd gnd cell_6t
Xbit_r66_c131 bl_131 br_131 wl_66 vdd gnd cell_6t
Xbit_r67_c131 bl_131 br_131 wl_67 vdd gnd cell_6t
Xbit_r68_c131 bl_131 br_131 wl_68 vdd gnd cell_6t
Xbit_r69_c131 bl_131 br_131 wl_69 vdd gnd cell_6t
Xbit_r70_c131 bl_131 br_131 wl_70 vdd gnd cell_6t
Xbit_r71_c131 bl_131 br_131 wl_71 vdd gnd cell_6t
Xbit_r72_c131 bl_131 br_131 wl_72 vdd gnd cell_6t
Xbit_r73_c131 bl_131 br_131 wl_73 vdd gnd cell_6t
Xbit_r74_c131 bl_131 br_131 wl_74 vdd gnd cell_6t
Xbit_r75_c131 bl_131 br_131 wl_75 vdd gnd cell_6t
Xbit_r76_c131 bl_131 br_131 wl_76 vdd gnd cell_6t
Xbit_r77_c131 bl_131 br_131 wl_77 vdd gnd cell_6t
Xbit_r78_c131 bl_131 br_131 wl_78 vdd gnd cell_6t
Xbit_r79_c131 bl_131 br_131 wl_79 vdd gnd cell_6t
Xbit_r80_c131 bl_131 br_131 wl_80 vdd gnd cell_6t
Xbit_r81_c131 bl_131 br_131 wl_81 vdd gnd cell_6t
Xbit_r82_c131 bl_131 br_131 wl_82 vdd gnd cell_6t
Xbit_r83_c131 bl_131 br_131 wl_83 vdd gnd cell_6t
Xbit_r84_c131 bl_131 br_131 wl_84 vdd gnd cell_6t
Xbit_r85_c131 bl_131 br_131 wl_85 vdd gnd cell_6t
Xbit_r86_c131 bl_131 br_131 wl_86 vdd gnd cell_6t
Xbit_r87_c131 bl_131 br_131 wl_87 vdd gnd cell_6t
Xbit_r88_c131 bl_131 br_131 wl_88 vdd gnd cell_6t
Xbit_r89_c131 bl_131 br_131 wl_89 vdd gnd cell_6t
Xbit_r90_c131 bl_131 br_131 wl_90 vdd gnd cell_6t
Xbit_r91_c131 bl_131 br_131 wl_91 vdd gnd cell_6t
Xbit_r92_c131 bl_131 br_131 wl_92 vdd gnd cell_6t
Xbit_r93_c131 bl_131 br_131 wl_93 vdd gnd cell_6t
Xbit_r94_c131 bl_131 br_131 wl_94 vdd gnd cell_6t
Xbit_r95_c131 bl_131 br_131 wl_95 vdd gnd cell_6t
Xbit_r96_c131 bl_131 br_131 wl_96 vdd gnd cell_6t
Xbit_r97_c131 bl_131 br_131 wl_97 vdd gnd cell_6t
Xbit_r98_c131 bl_131 br_131 wl_98 vdd gnd cell_6t
Xbit_r99_c131 bl_131 br_131 wl_99 vdd gnd cell_6t
Xbit_r100_c131 bl_131 br_131 wl_100 vdd gnd cell_6t
Xbit_r101_c131 bl_131 br_131 wl_101 vdd gnd cell_6t
Xbit_r102_c131 bl_131 br_131 wl_102 vdd gnd cell_6t
Xbit_r103_c131 bl_131 br_131 wl_103 vdd gnd cell_6t
Xbit_r104_c131 bl_131 br_131 wl_104 vdd gnd cell_6t
Xbit_r105_c131 bl_131 br_131 wl_105 vdd gnd cell_6t
Xbit_r106_c131 bl_131 br_131 wl_106 vdd gnd cell_6t
Xbit_r107_c131 bl_131 br_131 wl_107 vdd gnd cell_6t
Xbit_r108_c131 bl_131 br_131 wl_108 vdd gnd cell_6t
Xbit_r109_c131 bl_131 br_131 wl_109 vdd gnd cell_6t
Xbit_r110_c131 bl_131 br_131 wl_110 vdd gnd cell_6t
Xbit_r111_c131 bl_131 br_131 wl_111 vdd gnd cell_6t
Xbit_r112_c131 bl_131 br_131 wl_112 vdd gnd cell_6t
Xbit_r113_c131 bl_131 br_131 wl_113 vdd gnd cell_6t
Xbit_r114_c131 bl_131 br_131 wl_114 vdd gnd cell_6t
Xbit_r115_c131 bl_131 br_131 wl_115 vdd gnd cell_6t
Xbit_r116_c131 bl_131 br_131 wl_116 vdd gnd cell_6t
Xbit_r117_c131 bl_131 br_131 wl_117 vdd gnd cell_6t
Xbit_r118_c131 bl_131 br_131 wl_118 vdd gnd cell_6t
Xbit_r119_c131 bl_131 br_131 wl_119 vdd gnd cell_6t
Xbit_r120_c131 bl_131 br_131 wl_120 vdd gnd cell_6t
Xbit_r121_c131 bl_131 br_131 wl_121 vdd gnd cell_6t
Xbit_r122_c131 bl_131 br_131 wl_122 vdd gnd cell_6t
Xbit_r123_c131 bl_131 br_131 wl_123 vdd gnd cell_6t
Xbit_r124_c131 bl_131 br_131 wl_124 vdd gnd cell_6t
Xbit_r125_c131 bl_131 br_131 wl_125 vdd gnd cell_6t
Xbit_r126_c131 bl_131 br_131 wl_126 vdd gnd cell_6t
Xbit_r127_c131 bl_131 br_131 wl_127 vdd gnd cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd cell_6t
Xbit_r1_c132 bl_132 br_132 wl_1 vdd gnd cell_6t
Xbit_r2_c132 bl_132 br_132 wl_2 vdd gnd cell_6t
Xbit_r3_c132 bl_132 br_132 wl_3 vdd gnd cell_6t
Xbit_r4_c132 bl_132 br_132 wl_4 vdd gnd cell_6t
Xbit_r5_c132 bl_132 br_132 wl_5 vdd gnd cell_6t
Xbit_r6_c132 bl_132 br_132 wl_6 vdd gnd cell_6t
Xbit_r7_c132 bl_132 br_132 wl_7 vdd gnd cell_6t
Xbit_r8_c132 bl_132 br_132 wl_8 vdd gnd cell_6t
Xbit_r9_c132 bl_132 br_132 wl_9 vdd gnd cell_6t
Xbit_r10_c132 bl_132 br_132 wl_10 vdd gnd cell_6t
Xbit_r11_c132 bl_132 br_132 wl_11 vdd gnd cell_6t
Xbit_r12_c132 bl_132 br_132 wl_12 vdd gnd cell_6t
Xbit_r13_c132 bl_132 br_132 wl_13 vdd gnd cell_6t
Xbit_r14_c132 bl_132 br_132 wl_14 vdd gnd cell_6t
Xbit_r15_c132 bl_132 br_132 wl_15 vdd gnd cell_6t
Xbit_r16_c132 bl_132 br_132 wl_16 vdd gnd cell_6t
Xbit_r17_c132 bl_132 br_132 wl_17 vdd gnd cell_6t
Xbit_r18_c132 bl_132 br_132 wl_18 vdd gnd cell_6t
Xbit_r19_c132 bl_132 br_132 wl_19 vdd gnd cell_6t
Xbit_r20_c132 bl_132 br_132 wl_20 vdd gnd cell_6t
Xbit_r21_c132 bl_132 br_132 wl_21 vdd gnd cell_6t
Xbit_r22_c132 bl_132 br_132 wl_22 vdd gnd cell_6t
Xbit_r23_c132 bl_132 br_132 wl_23 vdd gnd cell_6t
Xbit_r24_c132 bl_132 br_132 wl_24 vdd gnd cell_6t
Xbit_r25_c132 bl_132 br_132 wl_25 vdd gnd cell_6t
Xbit_r26_c132 bl_132 br_132 wl_26 vdd gnd cell_6t
Xbit_r27_c132 bl_132 br_132 wl_27 vdd gnd cell_6t
Xbit_r28_c132 bl_132 br_132 wl_28 vdd gnd cell_6t
Xbit_r29_c132 bl_132 br_132 wl_29 vdd gnd cell_6t
Xbit_r30_c132 bl_132 br_132 wl_30 vdd gnd cell_6t
Xbit_r31_c132 bl_132 br_132 wl_31 vdd gnd cell_6t
Xbit_r32_c132 bl_132 br_132 wl_32 vdd gnd cell_6t
Xbit_r33_c132 bl_132 br_132 wl_33 vdd gnd cell_6t
Xbit_r34_c132 bl_132 br_132 wl_34 vdd gnd cell_6t
Xbit_r35_c132 bl_132 br_132 wl_35 vdd gnd cell_6t
Xbit_r36_c132 bl_132 br_132 wl_36 vdd gnd cell_6t
Xbit_r37_c132 bl_132 br_132 wl_37 vdd gnd cell_6t
Xbit_r38_c132 bl_132 br_132 wl_38 vdd gnd cell_6t
Xbit_r39_c132 bl_132 br_132 wl_39 vdd gnd cell_6t
Xbit_r40_c132 bl_132 br_132 wl_40 vdd gnd cell_6t
Xbit_r41_c132 bl_132 br_132 wl_41 vdd gnd cell_6t
Xbit_r42_c132 bl_132 br_132 wl_42 vdd gnd cell_6t
Xbit_r43_c132 bl_132 br_132 wl_43 vdd gnd cell_6t
Xbit_r44_c132 bl_132 br_132 wl_44 vdd gnd cell_6t
Xbit_r45_c132 bl_132 br_132 wl_45 vdd gnd cell_6t
Xbit_r46_c132 bl_132 br_132 wl_46 vdd gnd cell_6t
Xbit_r47_c132 bl_132 br_132 wl_47 vdd gnd cell_6t
Xbit_r48_c132 bl_132 br_132 wl_48 vdd gnd cell_6t
Xbit_r49_c132 bl_132 br_132 wl_49 vdd gnd cell_6t
Xbit_r50_c132 bl_132 br_132 wl_50 vdd gnd cell_6t
Xbit_r51_c132 bl_132 br_132 wl_51 vdd gnd cell_6t
Xbit_r52_c132 bl_132 br_132 wl_52 vdd gnd cell_6t
Xbit_r53_c132 bl_132 br_132 wl_53 vdd gnd cell_6t
Xbit_r54_c132 bl_132 br_132 wl_54 vdd gnd cell_6t
Xbit_r55_c132 bl_132 br_132 wl_55 vdd gnd cell_6t
Xbit_r56_c132 bl_132 br_132 wl_56 vdd gnd cell_6t
Xbit_r57_c132 bl_132 br_132 wl_57 vdd gnd cell_6t
Xbit_r58_c132 bl_132 br_132 wl_58 vdd gnd cell_6t
Xbit_r59_c132 bl_132 br_132 wl_59 vdd gnd cell_6t
Xbit_r60_c132 bl_132 br_132 wl_60 vdd gnd cell_6t
Xbit_r61_c132 bl_132 br_132 wl_61 vdd gnd cell_6t
Xbit_r62_c132 bl_132 br_132 wl_62 vdd gnd cell_6t
Xbit_r63_c132 bl_132 br_132 wl_63 vdd gnd cell_6t
Xbit_r64_c132 bl_132 br_132 wl_64 vdd gnd cell_6t
Xbit_r65_c132 bl_132 br_132 wl_65 vdd gnd cell_6t
Xbit_r66_c132 bl_132 br_132 wl_66 vdd gnd cell_6t
Xbit_r67_c132 bl_132 br_132 wl_67 vdd gnd cell_6t
Xbit_r68_c132 bl_132 br_132 wl_68 vdd gnd cell_6t
Xbit_r69_c132 bl_132 br_132 wl_69 vdd gnd cell_6t
Xbit_r70_c132 bl_132 br_132 wl_70 vdd gnd cell_6t
Xbit_r71_c132 bl_132 br_132 wl_71 vdd gnd cell_6t
Xbit_r72_c132 bl_132 br_132 wl_72 vdd gnd cell_6t
Xbit_r73_c132 bl_132 br_132 wl_73 vdd gnd cell_6t
Xbit_r74_c132 bl_132 br_132 wl_74 vdd gnd cell_6t
Xbit_r75_c132 bl_132 br_132 wl_75 vdd gnd cell_6t
Xbit_r76_c132 bl_132 br_132 wl_76 vdd gnd cell_6t
Xbit_r77_c132 bl_132 br_132 wl_77 vdd gnd cell_6t
Xbit_r78_c132 bl_132 br_132 wl_78 vdd gnd cell_6t
Xbit_r79_c132 bl_132 br_132 wl_79 vdd gnd cell_6t
Xbit_r80_c132 bl_132 br_132 wl_80 vdd gnd cell_6t
Xbit_r81_c132 bl_132 br_132 wl_81 vdd gnd cell_6t
Xbit_r82_c132 bl_132 br_132 wl_82 vdd gnd cell_6t
Xbit_r83_c132 bl_132 br_132 wl_83 vdd gnd cell_6t
Xbit_r84_c132 bl_132 br_132 wl_84 vdd gnd cell_6t
Xbit_r85_c132 bl_132 br_132 wl_85 vdd gnd cell_6t
Xbit_r86_c132 bl_132 br_132 wl_86 vdd gnd cell_6t
Xbit_r87_c132 bl_132 br_132 wl_87 vdd gnd cell_6t
Xbit_r88_c132 bl_132 br_132 wl_88 vdd gnd cell_6t
Xbit_r89_c132 bl_132 br_132 wl_89 vdd gnd cell_6t
Xbit_r90_c132 bl_132 br_132 wl_90 vdd gnd cell_6t
Xbit_r91_c132 bl_132 br_132 wl_91 vdd gnd cell_6t
Xbit_r92_c132 bl_132 br_132 wl_92 vdd gnd cell_6t
Xbit_r93_c132 bl_132 br_132 wl_93 vdd gnd cell_6t
Xbit_r94_c132 bl_132 br_132 wl_94 vdd gnd cell_6t
Xbit_r95_c132 bl_132 br_132 wl_95 vdd gnd cell_6t
Xbit_r96_c132 bl_132 br_132 wl_96 vdd gnd cell_6t
Xbit_r97_c132 bl_132 br_132 wl_97 vdd gnd cell_6t
Xbit_r98_c132 bl_132 br_132 wl_98 vdd gnd cell_6t
Xbit_r99_c132 bl_132 br_132 wl_99 vdd gnd cell_6t
Xbit_r100_c132 bl_132 br_132 wl_100 vdd gnd cell_6t
Xbit_r101_c132 bl_132 br_132 wl_101 vdd gnd cell_6t
Xbit_r102_c132 bl_132 br_132 wl_102 vdd gnd cell_6t
Xbit_r103_c132 bl_132 br_132 wl_103 vdd gnd cell_6t
Xbit_r104_c132 bl_132 br_132 wl_104 vdd gnd cell_6t
Xbit_r105_c132 bl_132 br_132 wl_105 vdd gnd cell_6t
Xbit_r106_c132 bl_132 br_132 wl_106 vdd gnd cell_6t
Xbit_r107_c132 bl_132 br_132 wl_107 vdd gnd cell_6t
Xbit_r108_c132 bl_132 br_132 wl_108 vdd gnd cell_6t
Xbit_r109_c132 bl_132 br_132 wl_109 vdd gnd cell_6t
Xbit_r110_c132 bl_132 br_132 wl_110 vdd gnd cell_6t
Xbit_r111_c132 bl_132 br_132 wl_111 vdd gnd cell_6t
Xbit_r112_c132 bl_132 br_132 wl_112 vdd gnd cell_6t
Xbit_r113_c132 bl_132 br_132 wl_113 vdd gnd cell_6t
Xbit_r114_c132 bl_132 br_132 wl_114 vdd gnd cell_6t
Xbit_r115_c132 bl_132 br_132 wl_115 vdd gnd cell_6t
Xbit_r116_c132 bl_132 br_132 wl_116 vdd gnd cell_6t
Xbit_r117_c132 bl_132 br_132 wl_117 vdd gnd cell_6t
Xbit_r118_c132 bl_132 br_132 wl_118 vdd gnd cell_6t
Xbit_r119_c132 bl_132 br_132 wl_119 vdd gnd cell_6t
Xbit_r120_c132 bl_132 br_132 wl_120 vdd gnd cell_6t
Xbit_r121_c132 bl_132 br_132 wl_121 vdd gnd cell_6t
Xbit_r122_c132 bl_132 br_132 wl_122 vdd gnd cell_6t
Xbit_r123_c132 bl_132 br_132 wl_123 vdd gnd cell_6t
Xbit_r124_c132 bl_132 br_132 wl_124 vdd gnd cell_6t
Xbit_r125_c132 bl_132 br_132 wl_125 vdd gnd cell_6t
Xbit_r126_c132 bl_132 br_132 wl_126 vdd gnd cell_6t
Xbit_r127_c132 bl_132 br_132 wl_127 vdd gnd cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd cell_6t
Xbit_r1_c133 bl_133 br_133 wl_1 vdd gnd cell_6t
Xbit_r2_c133 bl_133 br_133 wl_2 vdd gnd cell_6t
Xbit_r3_c133 bl_133 br_133 wl_3 vdd gnd cell_6t
Xbit_r4_c133 bl_133 br_133 wl_4 vdd gnd cell_6t
Xbit_r5_c133 bl_133 br_133 wl_5 vdd gnd cell_6t
Xbit_r6_c133 bl_133 br_133 wl_6 vdd gnd cell_6t
Xbit_r7_c133 bl_133 br_133 wl_7 vdd gnd cell_6t
Xbit_r8_c133 bl_133 br_133 wl_8 vdd gnd cell_6t
Xbit_r9_c133 bl_133 br_133 wl_9 vdd gnd cell_6t
Xbit_r10_c133 bl_133 br_133 wl_10 vdd gnd cell_6t
Xbit_r11_c133 bl_133 br_133 wl_11 vdd gnd cell_6t
Xbit_r12_c133 bl_133 br_133 wl_12 vdd gnd cell_6t
Xbit_r13_c133 bl_133 br_133 wl_13 vdd gnd cell_6t
Xbit_r14_c133 bl_133 br_133 wl_14 vdd gnd cell_6t
Xbit_r15_c133 bl_133 br_133 wl_15 vdd gnd cell_6t
Xbit_r16_c133 bl_133 br_133 wl_16 vdd gnd cell_6t
Xbit_r17_c133 bl_133 br_133 wl_17 vdd gnd cell_6t
Xbit_r18_c133 bl_133 br_133 wl_18 vdd gnd cell_6t
Xbit_r19_c133 bl_133 br_133 wl_19 vdd gnd cell_6t
Xbit_r20_c133 bl_133 br_133 wl_20 vdd gnd cell_6t
Xbit_r21_c133 bl_133 br_133 wl_21 vdd gnd cell_6t
Xbit_r22_c133 bl_133 br_133 wl_22 vdd gnd cell_6t
Xbit_r23_c133 bl_133 br_133 wl_23 vdd gnd cell_6t
Xbit_r24_c133 bl_133 br_133 wl_24 vdd gnd cell_6t
Xbit_r25_c133 bl_133 br_133 wl_25 vdd gnd cell_6t
Xbit_r26_c133 bl_133 br_133 wl_26 vdd gnd cell_6t
Xbit_r27_c133 bl_133 br_133 wl_27 vdd gnd cell_6t
Xbit_r28_c133 bl_133 br_133 wl_28 vdd gnd cell_6t
Xbit_r29_c133 bl_133 br_133 wl_29 vdd gnd cell_6t
Xbit_r30_c133 bl_133 br_133 wl_30 vdd gnd cell_6t
Xbit_r31_c133 bl_133 br_133 wl_31 vdd gnd cell_6t
Xbit_r32_c133 bl_133 br_133 wl_32 vdd gnd cell_6t
Xbit_r33_c133 bl_133 br_133 wl_33 vdd gnd cell_6t
Xbit_r34_c133 bl_133 br_133 wl_34 vdd gnd cell_6t
Xbit_r35_c133 bl_133 br_133 wl_35 vdd gnd cell_6t
Xbit_r36_c133 bl_133 br_133 wl_36 vdd gnd cell_6t
Xbit_r37_c133 bl_133 br_133 wl_37 vdd gnd cell_6t
Xbit_r38_c133 bl_133 br_133 wl_38 vdd gnd cell_6t
Xbit_r39_c133 bl_133 br_133 wl_39 vdd gnd cell_6t
Xbit_r40_c133 bl_133 br_133 wl_40 vdd gnd cell_6t
Xbit_r41_c133 bl_133 br_133 wl_41 vdd gnd cell_6t
Xbit_r42_c133 bl_133 br_133 wl_42 vdd gnd cell_6t
Xbit_r43_c133 bl_133 br_133 wl_43 vdd gnd cell_6t
Xbit_r44_c133 bl_133 br_133 wl_44 vdd gnd cell_6t
Xbit_r45_c133 bl_133 br_133 wl_45 vdd gnd cell_6t
Xbit_r46_c133 bl_133 br_133 wl_46 vdd gnd cell_6t
Xbit_r47_c133 bl_133 br_133 wl_47 vdd gnd cell_6t
Xbit_r48_c133 bl_133 br_133 wl_48 vdd gnd cell_6t
Xbit_r49_c133 bl_133 br_133 wl_49 vdd gnd cell_6t
Xbit_r50_c133 bl_133 br_133 wl_50 vdd gnd cell_6t
Xbit_r51_c133 bl_133 br_133 wl_51 vdd gnd cell_6t
Xbit_r52_c133 bl_133 br_133 wl_52 vdd gnd cell_6t
Xbit_r53_c133 bl_133 br_133 wl_53 vdd gnd cell_6t
Xbit_r54_c133 bl_133 br_133 wl_54 vdd gnd cell_6t
Xbit_r55_c133 bl_133 br_133 wl_55 vdd gnd cell_6t
Xbit_r56_c133 bl_133 br_133 wl_56 vdd gnd cell_6t
Xbit_r57_c133 bl_133 br_133 wl_57 vdd gnd cell_6t
Xbit_r58_c133 bl_133 br_133 wl_58 vdd gnd cell_6t
Xbit_r59_c133 bl_133 br_133 wl_59 vdd gnd cell_6t
Xbit_r60_c133 bl_133 br_133 wl_60 vdd gnd cell_6t
Xbit_r61_c133 bl_133 br_133 wl_61 vdd gnd cell_6t
Xbit_r62_c133 bl_133 br_133 wl_62 vdd gnd cell_6t
Xbit_r63_c133 bl_133 br_133 wl_63 vdd gnd cell_6t
Xbit_r64_c133 bl_133 br_133 wl_64 vdd gnd cell_6t
Xbit_r65_c133 bl_133 br_133 wl_65 vdd gnd cell_6t
Xbit_r66_c133 bl_133 br_133 wl_66 vdd gnd cell_6t
Xbit_r67_c133 bl_133 br_133 wl_67 vdd gnd cell_6t
Xbit_r68_c133 bl_133 br_133 wl_68 vdd gnd cell_6t
Xbit_r69_c133 bl_133 br_133 wl_69 vdd gnd cell_6t
Xbit_r70_c133 bl_133 br_133 wl_70 vdd gnd cell_6t
Xbit_r71_c133 bl_133 br_133 wl_71 vdd gnd cell_6t
Xbit_r72_c133 bl_133 br_133 wl_72 vdd gnd cell_6t
Xbit_r73_c133 bl_133 br_133 wl_73 vdd gnd cell_6t
Xbit_r74_c133 bl_133 br_133 wl_74 vdd gnd cell_6t
Xbit_r75_c133 bl_133 br_133 wl_75 vdd gnd cell_6t
Xbit_r76_c133 bl_133 br_133 wl_76 vdd gnd cell_6t
Xbit_r77_c133 bl_133 br_133 wl_77 vdd gnd cell_6t
Xbit_r78_c133 bl_133 br_133 wl_78 vdd gnd cell_6t
Xbit_r79_c133 bl_133 br_133 wl_79 vdd gnd cell_6t
Xbit_r80_c133 bl_133 br_133 wl_80 vdd gnd cell_6t
Xbit_r81_c133 bl_133 br_133 wl_81 vdd gnd cell_6t
Xbit_r82_c133 bl_133 br_133 wl_82 vdd gnd cell_6t
Xbit_r83_c133 bl_133 br_133 wl_83 vdd gnd cell_6t
Xbit_r84_c133 bl_133 br_133 wl_84 vdd gnd cell_6t
Xbit_r85_c133 bl_133 br_133 wl_85 vdd gnd cell_6t
Xbit_r86_c133 bl_133 br_133 wl_86 vdd gnd cell_6t
Xbit_r87_c133 bl_133 br_133 wl_87 vdd gnd cell_6t
Xbit_r88_c133 bl_133 br_133 wl_88 vdd gnd cell_6t
Xbit_r89_c133 bl_133 br_133 wl_89 vdd gnd cell_6t
Xbit_r90_c133 bl_133 br_133 wl_90 vdd gnd cell_6t
Xbit_r91_c133 bl_133 br_133 wl_91 vdd gnd cell_6t
Xbit_r92_c133 bl_133 br_133 wl_92 vdd gnd cell_6t
Xbit_r93_c133 bl_133 br_133 wl_93 vdd gnd cell_6t
Xbit_r94_c133 bl_133 br_133 wl_94 vdd gnd cell_6t
Xbit_r95_c133 bl_133 br_133 wl_95 vdd gnd cell_6t
Xbit_r96_c133 bl_133 br_133 wl_96 vdd gnd cell_6t
Xbit_r97_c133 bl_133 br_133 wl_97 vdd gnd cell_6t
Xbit_r98_c133 bl_133 br_133 wl_98 vdd gnd cell_6t
Xbit_r99_c133 bl_133 br_133 wl_99 vdd gnd cell_6t
Xbit_r100_c133 bl_133 br_133 wl_100 vdd gnd cell_6t
Xbit_r101_c133 bl_133 br_133 wl_101 vdd gnd cell_6t
Xbit_r102_c133 bl_133 br_133 wl_102 vdd gnd cell_6t
Xbit_r103_c133 bl_133 br_133 wl_103 vdd gnd cell_6t
Xbit_r104_c133 bl_133 br_133 wl_104 vdd gnd cell_6t
Xbit_r105_c133 bl_133 br_133 wl_105 vdd gnd cell_6t
Xbit_r106_c133 bl_133 br_133 wl_106 vdd gnd cell_6t
Xbit_r107_c133 bl_133 br_133 wl_107 vdd gnd cell_6t
Xbit_r108_c133 bl_133 br_133 wl_108 vdd gnd cell_6t
Xbit_r109_c133 bl_133 br_133 wl_109 vdd gnd cell_6t
Xbit_r110_c133 bl_133 br_133 wl_110 vdd gnd cell_6t
Xbit_r111_c133 bl_133 br_133 wl_111 vdd gnd cell_6t
Xbit_r112_c133 bl_133 br_133 wl_112 vdd gnd cell_6t
Xbit_r113_c133 bl_133 br_133 wl_113 vdd gnd cell_6t
Xbit_r114_c133 bl_133 br_133 wl_114 vdd gnd cell_6t
Xbit_r115_c133 bl_133 br_133 wl_115 vdd gnd cell_6t
Xbit_r116_c133 bl_133 br_133 wl_116 vdd gnd cell_6t
Xbit_r117_c133 bl_133 br_133 wl_117 vdd gnd cell_6t
Xbit_r118_c133 bl_133 br_133 wl_118 vdd gnd cell_6t
Xbit_r119_c133 bl_133 br_133 wl_119 vdd gnd cell_6t
Xbit_r120_c133 bl_133 br_133 wl_120 vdd gnd cell_6t
Xbit_r121_c133 bl_133 br_133 wl_121 vdd gnd cell_6t
Xbit_r122_c133 bl_133 br_133 wl_122 vdd gnd cell_6t
Xbit_r123_c133 bl_133 br_133 wl_123 vdd gnd cell_6t
Xbit_r124_c133 bl_133 br_133 wl_124 vdd gnd cell_6t
Xbit_r125_c133 bl_133 br_133 wl_125 vdd gnd cell_6t
Xbit_r126_c133 bl_133 br_133 wl_126 vdd gnd cell_6t
Xbit_r127_c133 bl_133 br_133 wl_127 vdd gnd cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd cell_6t
Xbit_r1_c134 bl_134 br_134 wl_1 vdd gnd cell_6t
Xbit_r2_c134 bl_134 br_134 wl_2 vdd gnd cell_6t
Xbit_r3_c134 bl_134 br_134 wl_3 vdd gnd cell_6t
Xbit_r4_c134 bl_134 br_134 wl_4 vdd gnd cell_6t
Xbit_r5_c134 bl_134 br_134 wl_5 vdd gnd cell_6t
Xbit_r6_c134 bl_134 br_134 wl_6 vdd gnd cell_6t
Xbit_r7_c134 bl_134 br_134 wl_7 vdd gnd cell_6t
Xbit_r8_c134 bl_134 br_134 wl_8 vdd gnd cell_6t
Xbit_r9_c134 bl_134 br_134 wl_9 vdd gnd cell_6t
Xbit_r10_c134 bl_134 br_134 wl_10 vdd gnd cell_6t
Xbit_r11_c134 bl_134 br_134 wl_11 vdd gnd cell_6t
Xbit_r12_c134 bl_134 br_134 wl_12 vdd gnd cell_6t
Xbit_r13_c134 bl_134 br_134 wl_13 vdd gnd cell_6t
Xbit_r14_c134 bl_134 br_134 wl_14 vdd gnd cell_6t
Xbit_r15_c134 bl_134 br_134 wl_15 vdd gnd cell_6t
Xbit_r16_c134 bl_134 br_134 wl_16 vdd gnd cell_6t
Xbit_r17_c134 bl_134 br_134 wl_17 vdd gnd cell_6t
Xbit_r18_c134 bl_134 br_134 wl_18 vdd gnd cell_6t
Xbit_r19_c134 bl_134 br_134 wl_19 vdd gnd cell_6t
Xbit_r20_c134 bl_134 br_134 wl_20 vdd gnd cell_6t
Xbit_r21_c134 bl_134 br_134 wl_21 vdd gnd cell_6t
Xbit_r22_c134 bl_134 br_134 wl_22 vdd gnd cell_6t
Xbit_r23_c134 bl_134 br_134 wl_23 vdd gnd cell_6t
Xbit_r24_c134 bl_134 br_134 wl_24 vdd gnd cell_6t
Xbit_r25_c134 bl_134 br_134 wl_25 vdd gnd cell_6t
Xbit_r26_c134 bl_134 br_134 wl_26 vdd gnd cell_6t
Xbit_r27_c134 bl_134 br_134 wl_27 vdd gnd cell_6t
Xbit_r28_c134 bl_134 br_134 wl_28 vdd gnd cell_6t
Xbit_r29_c134 bl_134 br_134 wl_29 vdd gnd cell_6t
Xbit_r30_c134 bl_134 br_134 wl_30 vdd gnd cell_6t
Xbit_r31_c134 bl_134 br_134 wl_31 vdd gnd cell_6t
Xbit_r32_c134 bl_134 br_134 wl_32 vdd gnd cell_6t
Xbit_r33_c134 bl_134 br_134 wl_33 vdd gnd cell_6t
Xbit_r34_c134 bl_134 br_134 wl_34 vdd gnd cell_6t
Xbit_r35_c134 bl_134 br_134 wl_35 vdd gnd cell_6t
Xbit_r36_c134 bl_134 br_134 wl_36 vdd gnd cell_6t
Xbit_r37_c134 bl_134 br_134 wl_37 vdd gnd cell_6t
Xbit_r38_c134 bl_134 br_134 wl_38 vdd gnd cell_6t
Xbit_r39_c134 bl_134 br_134 wl_39 vdd gnd cell_6t
Xbit_r40_c134 bl_134 br_134 wl_40 vdd gnd cell_6t
Xbit_r41_c134 bl_134 br_134 wl_41 vdd gnd cell_6t
Xbit_r42_c134 bl_134 br_134 wl_42 vdd gnd cell_6t
Xbit_r43_c134 bl_134 br_134 wl_43 vdd gnd cell_6t
Xbit_r44_c134 bl_134 br_134 wl_44 vdd gnd cell_6t
Xbit_r45_c134 bl_134 br_134 wl_45 vdd gnd cell_6t
Xbit_r46_c134 bl_134 br_134 wl_46 vdd gnd cell_6t
Xbit_r47_c134 bl_134 br_134 wl_47 vdd gnd cell_6t
Xbit_r48_c134 bl_134 br_134 wl_48 vdd gnd cell_6t
Xbit_r49_c134 bl_134 br_134 wl_49 vdd gnd cell_6t
Xbit_r50_c134 bl_134 br_134 wl_50 vdd gnd cell_6t
Xbit_r51_c134 bl_134 br_134 wl_51 vdd gnd cell_6t
Xbit_r52_c134 bl_134 br_134 wl_52 vdd gnd cell_6t
Xbit_r53_c134 bl_134 br_134 wl_53 vdd gnd cell_6t
Xbit_r54_c134 bl_134 br_134 wl_54 vdd gnd cell_6t
Xbit_r55_c134 bl_134 br_134 wl_55 vdd gnd cell_6t
Xbit_r56_c134 bl_134 br_134 wl_56 vdd gnd cell_6t
Xbit_r57_c134 bl_134 br_134 wl_57 vdd gnd cell_6t
Xbit_r58_c134 bl_134 br_134 wl_58 vdd gnd cell_6t
Xbit_r59_c134 bl_134 br_134 wl_59 vdd gnd cell_6t
Xbit_r60_c134 bl_134 br_134 wl_60 vdd gnd cell_6t
Xbit_r61_c134 bl_134 br_134 wl_61 vdd gnd cell_6t
Xbit_r62_c134 bl_134 br_134 wl_62 vdd gnd cell_6t
Xbit_r63_c134 bl_134 br_134 wl_63 vdd gnd cell_6t
Xbit_r64_c134 bl_134 br_134 wl_64 vdd gnd cell_6t
Xbit_r65_c134 bl_134 br_134 wl_65 vdd gnd cell_6t
Xbit_r66_c134 bl_134 br_134 wl_66 vdd gnd cell_6t
Xbit_r67_c134 bl_134 br_134 wl_67 vdd gnd cell_6t
Xbit_r68_c134 bl_134 br_134 wl_68 vdd gnd cell_6t
Xbit_r69_c134 bl_134 br_134 wl_69 vdd gnd cell_6t
Xbit_r70_c134 bl_134 br_134 wl_70 vdd gnd cell_6t
Xbit_r71_c134 bl_134 br_134 wl_71 vdd gnd cell_6t
Xbit_r72_c134 bl_134 br_134 wl_72 vdd gnd cell_6t
Xbit_r73_c134 bl_134 br_134 wl_73 vdd gnd cell_6t
Xbit_r74_c134 bl_134 br_134 wl_74 vdd gnd cell_6t
Xbit_r75_c134 bl_134 br_134 wl_75 vdd gnd cell_6t
Xbit_r76_c134 bl_134 br_134 wl_76 vdd gnd cell_6t
Xbit_r77_c134 bl_134 br_134 wl_77 vdd gnd cell_6t
Xbit_r78_c134 bl_134 br_134 wl_78 vdd gnd cell_6t
Xbit_r79_c134 bl_134 br_134 wl_79 vdd gnd cell_6t
Xbit_r80_c134 bl_134 br_134 wl_80 vdd gnd cell_6t
Xbit_r81_c134 bl_134 br_134 wl_81 vdd gnd cell_6t
Xbit_r82_c134 bl_134 br_134 wl_82 vdd gnd cell_6t
Xbit_r83_c134 bl_134 br_134 wl_83 vdd gnd cell_6t
Xbit_r84_c134 bl_134 br_134 wl_84 vdd gnd cell_6t
Xbit_r85_c134 bl_134 br_134 wl_85 vdd gnd cell_6t
Xbit_r86_c134 bl_134 br_134 wl_86 vdd gnd cell_6t
Xbit_r87_c134 bl_134 br_134 wl_87 vdd gnd cell_6t
Xbit_r88_c134 bl_134 br_134 wl_88 vdd gnd cell_6t
Xbit_r89_c134 bl_134 br_134 wl_89 vdd gnd cell_6t
Xbit_r90_c134 bl_134 br_134 wl_90 vdd gnd cell_6t
Xbit_r91_c134 bl_134 br_134 wl_91 vdd gnd cell_6t
Xbit_r92_c134 bl_134 br_134 wl_92 vdd gnd cell_6t
Xbit_r93_c134 bl_134 br_134 wl_93 vdd gnd cell_6t
Xbit_r94_c134 bl_134 br_134 wl_94 vdd gnd cell_6t
Xbit_r95_c134 bl_134 br_134 wl_95 vdd gnd cell_6t
Xbit_r96_c134 bl_134 br_134 wl_96 vdd gnd cell_6t
Xbit_r97_c134 bl_134 br_134 wl_97 vdd gnd cell_6t
Xbit_r98_c134 bl_134 br_134 wl_98 vdd gnd cell_6t
Xbit_r99_c134 bl_134 br_134 wl_99 vdd gnd cell_6t
Xbit_r100_c134 bl_134 br_134 wl_100 vdd gnd cell_6t
Xbit_r101_c134 bl_134 br_134 wl_101 vdd gnd cell_6t
Xbit_r102_c134 bl_134 br_134 wl_102 vdd gnd cell_6t
Xbit_r103_c134 bl_134 br_134 wl_103 vdd gnd cell_6t
Xbit_r104_c134 bl_134 br_134 wl_104 vdd gnd cell_6t
Xbit_r105_c134 bl_134 br_134 wl_105 vdd gnd cell_6t
Xbit_r106_c134 bl_134 br_134 wl_106 vdd gnd cell_6t
Xbit_r107_c134 bl_134 br_134 wl_107 vdd gnd cell_6t
Xbit_r108_c134 bl_134 br_134 wl_108 vdd gnd cell_6t
Xbit_r109_c134 bl_134 br_134 wl_109 vdd gnd cell_6t
Xbit_r110_c134 bl_134 br_134 wl_110 vdd gnd cell_6t
Xbit_r111_c134 bl_134 br_134 wl_111 vdd gnd cell_6t
Xbit_r112_c134 bl_134 br_134 wl_112 vdd gnd cell_6t
Xbit_r113_c134 bl_134 br_134 wl_113 vdd gnd cell_6t
Xbit_r114_c134 bl_134 br_134 wl_114 vdd gnd cell_6t
Xbit_r115_c134 bl_134 br_134 wl_115 vdd gnd cell_6t
Xbit_r116_c134 bl_134 br_134 wl_116 vdd gnd cell_6t
Xbit_r117_c134 bl_134 br_134 wl_117 vdd gnd cell_6t
Xbit_r118_c134 bl_134 br_134 wl_118 vdd gnd cell_6t
Xbit_r119_c134 bl_134 br_134 wl_119 vdd gnd cell_6t
Xbit_r120_c134 bl_134 br_134 wl_120 vdd gnd cell_6t
Xbit_r121_c134 bl_134 br_134 wl_121 vdd gnd cell_6t
Xbit_r122_c134 bl_134 br_134 wl_122 vdd gnd cell_6t
Xbit_r123_c134 bl_134 br_134 wl_123 vdd gnd cell_6t
Xbit_r124_c134 bl_134 br_134 wl_124 vdd gnd cell_6t
Xbit_r125_c134 bl_134 br_134 wl_125 vdd gnd cell_6t
Xbit_r126_c134 bl_134 br_134 wl_126 vdd gnd cell_6t
Xbit_r127_c134 bl_134 br_134 wl_127 vdd gnd cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd cell_6t
Xbit_r1_c135 bl_135 br_135 wl_1 vdd gnd cell_6t
Xbit_r2_c135 bl_135 br_135 wl_2 vdd gnd cell_6t
Xbit_r3_c135 bl_135 br_135 wl_3 vdd gnd cell_6t
Xbit_r4_c135 bl_135 br_135 wl_4 vdd gnd cell_6t
Xbit_r5_c135 bl_135 br_135 wl_5 vdd gnd cell_6t
Xbit_r6_c135 bl_135 br_135 wl_6 vdd gnd cell_6t
Xbit_r7_c135 bl_135 br_135 wl_7 vdd gnd cell_6t
Xbit_r8_c135 bl_135 br_135 wl_8 vdd gnd cell_6t
Xbit_r9_c135 bl_135 br_135 wl_9 vdd gnd cell_6t
Xbit_r10_c135 bl_135 br_135 wl_10 vdd gnd cell_6t
Xbit_r11_c135 bl_135 br_135 wl_11 vdd gnd cell_6t
Xbit_r12_c135 bl_135 br_135 wl_12 vdd gnd cell_6t
Xbit_r13_c135 bl_135 br_135 wl_13 vdd gnd cell_6t
Xbit_r14_c135 bl_135 br_135 wl_14 vdd gnd cell_6t
Xbit_r15_c135 bl_135 br_135 wl_15 vdd gnd cell_6t
Xbit_r16_c135 bl_135 br_135 wl_16 vdd gnd cell_6t
Xbit_r17_c135 bl_135 br_135 wl_17 vdd gnd cell_6t
Xbit_r18_c135 bl_135 br_135 wl_18 vdd gnd cell_6t
Xbit_r19_c135 bl_135 br_135 wl_19 vdd gnd cell_6t
Xbit_r20_c135 bl_135 br_135 wl_20 vdd gnd cell_6t
Xbit_r21_c135 bl_135 br_135 wl_21 vdd gnd cell_6t
Xbit_r22_c135 bl_135 br_135 wl_22 vdd gnd cell_6t
Xbit_r23_c135 bl_135 br_135 wl_23 vdd gnd cell_6t
Xbit_r24_c135 bl_135 br_135 wl_24 vdd gnd cell_6t
Xbit_r25_c135 bl_135 br_135 wl_25 vdd gnd cell_6t
Xbit_r26_c135 bl_135 br_135 wl_26 vdd gnd cell_6t
Xbit_r27_c135 bl_135 br_135 wl_27 vdd gnd cell_6t
Xbit_r28_c135 bl_135 br_135 wl_28 vdd gnd cell_6t
Xbit_r29_c135 bl_135 br_135 wl_29 vdd gnd cell_6t
Xbit_r30_c135 bl_135 br_135 wl_30 vdd gnd cell_6t
Xbit_r31_c135 bl_135 br_135 wl_31 vdd gnd cell_6t
Xbit_r32_c135 bl_135 br_135 wl_32 vdd gnd cell_6t
Xbit_r33_c135 bl_135 br_135 wl_33 vdd gnd cell_6t
Xbit_r34_c135 bl_135 br_135 wl_34 vdd gnd cell_6t
Xbit_r35_c135 bl_135 br_135 wl_35 vdd gnd cell_6t
Xbit_r36_c135 bl_135 br_135 wl_36 vdd gnd cell_6t
Xbit_r37_c135 bl_135 br_135 wl_37 vdd gnd cell_6t
Xbit_r38_c135 bl_135 br_135 wl_38 vdd gnd cell_6t
Xbit_r39_c135 bl_135 br_135 wl_39 vdd gnd cell_6t
Xbit_r40_c135 bl_135 br_135 wl_40 vdd gnd cell_6t
Xbit_r41_c135 bl_135 br_135 wl_41 vdd gnd cell_6t
Xbit_r42_c135 bl_135 br_135 wl_42 vdd gnd cell_6t
Xbit_r43_c135 bl_135 br_135 wl_43 vdd gnd cell_6t
Xbit_r44_c135 bl_135 br_135 wl_44 vdd gnd cell_6t
Xbit_r45_c135 bl_135 br_135 wl_45 vdd gnd cell_6t
Xbit_r46_c135 bl_135 br_135 wl_46 vdd gnd cell_6t
Xbit_r47_c135 bl_135 br_135 wl_47 vdd gnd cell_6t
Xbit_r48_c135 bl_135 br_135 wl_48 vdd gnd cell_6t
Xbit_r49_c135 bl_135 br_135 wl_49 vdd gnd cell_6t
Xbit_r50_c135 bl_135 br_135 wl_50 vdd gnd cell_6t
Xbit_r51_c135 bl_135 br_135 wl_51 vdd gnd cell_6t
Xbit_r52_c135 bl_135 br_135 wl_52 vdd gnd cell_6t
Xbit_r53_c135 bl_135 br_135 wl_53 vdd gnd cell_6t
Xbit_r54_c135 bl_135 br_135 wl_54 vdd gnd cell_6t
Xbit_r55_c135 bl_135 br_135 wl_55 vdd gnd cell_6t
Xbit_r56_c135 bl_135 br_135 wl_56 vdd gnd cell_6t
Xbit_r57_c135 bl_135 br_135 wl_57 vdd gnd cell_6t
Xbit_r58_c135 bl_135 br_135 wl_58 vdd gnd cell_6t
Xbit_r59_c135 bl_135 br_135 wl_59 vdd gnd cell_6t
Xbit_r60_c135 bl_135 br_135 wl_60 vdd gnd cell_6t
Xbit_r61_c135 bl_135 br_135 wl_61 vdd gnd cell_6t
Xbit_r62_c135 bl_135 br_135 wl_62 vdd gnd cell_6t
Xbit_r63_c135 bl_135 br_135 wl_63 vdd gnd cell_6t
Xbit_r64_c135 bl_135 br_135 wl_64 vdd gnd cell_6t
Xbit_r65_c135 bl_135 br_135 wl_65 vdd gnd cell_6t
Xbit_r66_c135 bl_135 br_135 wl_66 vdd gnd cell_6t
Xbit_r67_c135 bl_135 br_135 wl_67 vdd gnd cell_6t
Xbit_r68_c135 bl_135 br_135 wl_68 vdd gnd cell_6t
Xbit_r69_c135 bl_135 br_135 wl_69 vdd gnd cell_6t
Xbit_r70_c135 bl_135 br_135 wl_70 vdd gnd cell_6t
Xbit_r71_c135 bl_135 br_135 wl_71 vdd gnd cell_6t
Xbit_r72_c135 bl_135 br_135 wl_72 vdd gnd cell_6t
Xbit_r73_c135 bl_135 br_135 wl_73 vdd gnd cell_6t
Xbit_r74_c135 bl_135 br_135 wl_74 vdd gnd cell_6t
Xbit_r75_c135 bl_135 br_135 wl_75 vdd gnd cell_6t
Xbit_r76_c135 bl_135 br_135 wl_76 vdd gnd cell_6t
Xbit_r77_c135 bl_135 br_135 wl_77 vdd gnd cell_6t
Xbit_r78_c135 bl_135 br_135 wl_78 vdd gnd cell_6t
Xbit_r79_c135 bl_135 br_135 wl_79 vdd gnd cell_6t
Xbit_r80_c135 bl_135 br_135 wl_80 vdd gnd cell_6t
Xbit_r81_c135 bl_135 br_135 wl_81 vdd gnd cell_6t
Xbit_r82_c135 bl_135 br_135 wl_82 vdd gnd cell_6t
Xbit_r83_c135 bl_135 br_135 wl_83 vdd gnd cell_6t
Xbit_r84_c135 bl_135 br_135 wl_84 vdd gnd cell_6t
Xbit_r85_c135 bl_135 br_135 wl_85 vdd gnd cell_6t
Xbit_r86_c135 bl_135 br_135 wl_86 vdd gnd cell_6t
Xbit_r87_c135 bl_135 br_135 wl_87 vdd gnd cell_6t
Xbit_r88_c135 bl_135 br_135 wl_88 vdd gnd cell_6t
Xbit_r89_c135 bl_135 br_135 wl_89 vdd gnd cell_6t
Xbit_r90_c135 bl_135 br_135 wl_90 vdd gnd cell_6t
Xbit_r91_c135 bl_135 br_135 wl_91 vdd gnd cell_6t
Xbit_r92_c135 bl_135 br_135 wl_92 vdd gnd cell_6t
Xbit_r93_c135 bl_135 br_135 wl_93 vdd gnd cell_6t
Xbit_r94_c135 bl_135 br_135 wl_94 vdd gnd cell_6t
Xbit_r95_c135 bl_135 br_135 wl_95 vdd gnd cell_6t
Xbit_r96_c135 bl_135 br_135 wl_96 vdd gnd cell_6t
Xbit_r97_c135 bl_135 br_135 wl_97 vdd gnd cell_6t
Xbit_r98_c135 bl_135 br_135 wl_98 vdd gnd cell_6t
Xbit_r99_c135 bl_135 br_135 wl_99 vdd gnd cell_6t
Xbit_r100_c135 bl_135 br_135 wl_100 vdd gnd cell_6t
Xbit_r101_c135 bl_135 br_135 wl_101 vdd gnd cell_6t
Xbit_r102_c135 bl_135 br_135 wl_102 vdd gnd cell_6t
Xbit_r103_c135 bl_135 br_135 wl_103 vdd gnd cell_6t
Xbit_r104_c135 bl_135 br_135 wl_104 vdd gnd cell_6t
Xbit_r105_c135 bl_135 br_135 wl_105 vdd gnd cell_6t
Xbit_r106_c135 bl_135 br_135 wl_106 vdd gnd cell_6t
Xbit_r107_c135 bl_135 br_135 wl_107 vdd gnd cell_6t
Xbit_r108_c135 bl_135 br_135 wl_108 vdd gnd cell_6t
Xbit_r109_c135 bl_135 br_135 wl_109 vdd gnd cell_6t
Xbit_r110_c135 bl_135 br_135 wl_110 vdd gnd cell_6t
Xbit_r111_c135 bl_135 br_135 wl_111 vdd gnd cell_6t
Xbit_r112_c135 bl_135 br_135 wl_112 vdd gnd cell_6t
Xbit_r113_c135 bl_135 br_135 wl_113 vdd gnd cell_6t
Xbit_r114_c135 bl_135 br_135 wl_114 vdd gnd cell_6t
Xbit_r115_c135 bl_135 br_135 wl_115 vdd gnd cell_6t
Xbit_r116_c135 bl_135 br_135 wl_116 vdd gnd cell_6t
Xbit_r117_c135 bl_135 br_135 wl_117 vdd gnd cell_6t
Xbit_r118_c135 bl_135 br_135 wl_118 vdd gnd cell_6t
Xbit_r119_c135 bl_135 br_135 wl_119 vdd gnd cell_6t
Xbit_r120_c135 bl_135 br_135 wl_120 vdd gnd cell_6t
Xbit_r121_c135 bl_135 br_135 wl_121 vdd gnd cell_6t
Xbit_r122_c135 bl_135 br_135 wl_122 vdd gnd cell_6t
Xbit_r123_c135 bl_135 br_135 wl_123 vdd gnd cell_6t
Xbit_r124_c135 bl_135 br_135 wl_124 vdd gnd cell_6t
Xbit_r125_c135 bl_135 br_135 wl_125 vdd gnd cell_6t
Xbit_r126_c135 bl_135 br_135 wl_126 vdd gnd cell_6t
Xbit_r127_c135 bl_135 br_135 wl_127 vdd gnd cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd cell_6t
Xbit_r1_c136 bl_136 br_136 wl_1 vdd gnd cell_6t
Xbit_r2_c136 bl_136 br_136 wl_2 vdd gnd cell_6t
Xbit_r3_c136 bl_136 br_136 wl_3 vdd gnd cell_6t
Xbit_r4_c136 bl_136 br_136 wl_4 vdd gnd cell_6t
Xbit_r5_c136 bl_136 br_136 wl_5 vdd gnd cell_6t
Xbit_r6_c136 bl_136 br_136 wl_6 vdd gnd cell_6t
Xbit_r7_c136 bl_136 br_136 wl_7 vdd gnd cell_6t
Xbit_r8_c136 bl_136 br_136 wl_8 vdd gnd cell_6t
Xbit_r9_c136 bl_136 br_136 wl_9 vdd gnd cell_6t
Xbit_r10_c136 bl_136 br_136 wl_10 vdd gnd cell_6t
Xbit_r11_c136 bl_136 br_136 wl_11 vdd gnd cell_6t
Xbit_r12_c136 bl_136 br_136 wl_12 vdd gnd cell_6t
Xbit_r13_c136 bl_136 br_136 wl_13 vdd gnd cell_6t
Xbit_r14_c136 bl_136 br_136 wl_14 vdd gnd cell_6t
Xbit_r15_c136 bl_136 br_136 wl_15 vdd gnd cell_6t
Xbit_r16_c136 bl_136 br_136 wl_16 vdd gnd cell_6t
Xbit_r17_c136 bl_136 br_136 wl_17 vdd gnd cell_6t
Xbit_r18_c136 bl_136 br_136 wl_18 vdd gnd cell_6t
Xbit_r19_c136 bl_136 br_136 wl_19 vdd gnd cell_6t
Xbit_r20_c136 bl_136 br_136 wl_20 vdd gnd cell_6t
Xbit_r21_c136 bl_136 br_136 wl_21 vdd gnd cell_6t
Xbit_r22_c136 bl_136 br_136 wl_22 vdd gnd cell_6t
Xbit_r23_c136 bl_136 br_136 wl_23 vdd gnd cell_6t
Xbit_r24_c136 bl_136 br_136 wl_24 vdd gnd cell_6t
Xbit_r25_c136 bl_136 br_136 wl_25 vdd gnd cell_6t
Xbit_r26_c136 bl_136 br_136 wl_26 vdd gnd cell_6t
Xbit_r27_c136 bl_136 br_136 wl_27 vdd gnd cell_6t
Xbit_r28_c136 bl_136 br_136 wl_28 vdd gnd cell_6t
Xbit_r29_c136 bl_136 br_136 wl_29 vdd gnd cell_6t
Xbit_r30_c136 bl_136 br_136 wl_30 vdd gnd cell_6t
Xbit_r31_c136 bl_136 br_136 wl_31 vdd gnd cell_6t
Xbit_r32_c136 bl_136 br_136 wl_32 vdd gnd cell_6t
Xbit_r33_c136 bl_136 br_136 wl_33 vdd gnd cell_6t
Xbit_r34_c136 bl_136 br_136 wl_34 vdd gnd cell_6t
Xbit_r35_c136 bl_136 br_136 wl_35 vdd gnd cell_6t
Xbit_r36_c136 bl_136 br_136 wl_36 vdd gnd cell_6t
Xbit_r37_c136 bl_136 br_136 wl_37 vdd gnd cell_6t
Xbit_r38_c136 bl_136 br_136 wl_38 vdd gnd cell_6t
Xbit_r39_c136 bl_136 br_136 wl_39 vdd gnd cell_6t
Xbit_r40_c136 bl_136 br_136 wl_40 vdd gnd cell_6t
Xbit_r41_c136 bl_136 br_136 wl_41 vdd gnd cell_6t
Xbit_r42_c136 bl_136 br_136 wl_42 vdd gnd cell_6t
Xbit_r43_c136 bl_136 br_136 wl_43 vdd gnd cell_6t
Xbit_r44_c136 bl_136 br_136 wl_44 vdd gnd cell_6t
Xbit_r45_c136 bl_136 br_136 wl_45 vdd gnd cell_6t
Xbit_r46_c136 bl_136 br_136 wl_46 vdd gnd cell_6t
Xbit_r47_c136 bl_136 br_136 wl_47 vdd gnd cell_6t
Xbit_r48_c136 bl_136 br_136 wl_48 vdd gnd cell_6t
Xbit_r49_c136 bl_136 br_136 wl_49 vdd gnd cell_6t
Xbit_r50_c136 bl_136 br_136 wl_50 vdd gnd cell_6t
Xbit_r51_c136 bl_136 br_136 wl_51 vdd gnd cell_6t
Xbit_r52_c136 bl_136 br_136 wl_52 vdd gnd cell_6t
Xbit_r53_c136 bl_136 br_136 wl_53 vdd gnd cell_6t
Xbit_r54_c136 bl_136 br_136 wl_54 vdd gnd cell_6t
Xbit_r55_c136 bl_136 br_136 wl_55 vdd gnd cell_6t
Xbit_r56_c136 bl_136 br_136 wl_56 vdd gnd cell_6t
Xbit_r57_c136 bl_136 br_136 wl_57 vdd gnd cell_6t
Xbit_r58_c136 bl_136 br_136 wl_58 vdd gnd cell_6t
Xbit_r59_c136 bl_136 br_136 wl_59 vdd gnd cell_6t
Xbit_r60_c136 bl_136 br_136 wl_60 vdd gnd cell_6t
Xbit_r61_c136 bl_136 br_136 wl_61 vdd gnd cell_6t
Xbit_r62_c136 bl_136 br_136 wl_62 vdd gnd cell_6t
Xbit_r63_c136 bl_136 br_136 wl_63 vdd gnd cell_6t
Xbit_r64_c136 bl_136 br_136 wl_64 vdd gnd cell_6t
Xbit_r65_c136 bl_136 br_136 wl_65 vdd gnd cell_6t
Xbit_r66_c136 bl_136 br_136 wl_66 vdd gnd cell_6t
Xbit_r67_c136 bl_136 br_136 wl_67 vdd gnd cell_6t
Xbit_r68_c136 bl_136 br_136 wl_68 vdd gnd cell_6t
Xbit_r69_c136 bl_136 br_136 wl_69 vdd gnd cell_6t
Xbit_r70_c136 bl_136 br_136 wl_70 vdd gnd cell_6t
Xbit_r71_c136 bl_136 br_136 wl_71 vdd gnd cell_6t
Xbit_r72_c136 bl_136 br_136 wl_72 vdd gnd cell_6t
Xbit_r73_c136 bl_136 br_136 wl_73 vdd gnd cell_6t
Xbit_r74_c136 bl_136 br_136 wl_74 vdd gnd cell_6t
Xbit_r75_c136 bl_136 br_136 wl_75 vdd gnd cell_6t
Xbit_r76_c136 bl_136 br_136 wl_76 vdd gnd cell_6t
Xbit_r77_c136 bl_136 br_136 wl_77 vdd gnd cell_6t
Xbit_r78_c136 bl_136 br_136 wl_78 vdd gnd cell_6t
Xbit_r79_c136 bl_136 br_136 wl_79 vdd gnd cell_6t
Xbit_r80_c136 bl_136 br_136 wl_80 vdd gnd cell_6t
Xbit_r81_c136 bl_136 br_136 wl_81 vdd gnd cell_6t
Xbit_r82_c136 bl_136 br_136 wl_82 vdd gnd cell_6t
Xbit_r83_c136 bl_136 br_136 wl_83 vdd gnd cell_6t
Xbit_r84_c136 bl_136 br_136 wl_84 vdd gnd cell_6t
Xbit_r85_c136 bl_136 br_136 wl_85 vdd gnd cell_6t
Xbit_r86_c136 bl_136 br_136 wl_86 vdd gnd cell_6t
Xbit_r87_c136 bl_136 br_136 wl_87 vdd gnd cell_6t
Xbit_r88_c136 bl_136 br_136 wl_88 vdd gnd cell_6t
Xbit_r89_c136 bl_136 br_136 wl_89 vdd gnd cell_6t
Xbit_r90_c136 bl_136 br_136 wl_90 vdd gnd cell_6t
Xbit_r91_c136 bl_136 br_136 wl_91 vdd gnd cell_6t
Xbit_r92_c136 bl_136 br_136 wl_92 vdd gnd cell_6t
Xbit_r93_c136 bl_136 br_136 wl_93 vdd gnd cell_6t
Xbit_r94_c136 bl_136 br_136 wl_94 vdd gnd cell_6t
Xbit_r95_c136 bl_136 br_136 wl_95 vdd gnd cell_6t
Xbit_r96_c136 bl_136 br_136 wl_96 vdd gnd cell_6t
Xbit_r97_c136 bl_136 br_136 wl_97 vdd gnd cell_6t
Xbit_r98_c136 bl_136 br_136 wl_98 vdd gnd cell_6t
Xbit_r99_c136 bl_136 br_136 wl_99 vdd gnd cell_6t
Xbit_r100_c136 bl_136 br_136 wl_100 vdd gnd cell_6t
Xbit_r101_c136 bl_136 br_136 wl_101 vdd gnd cell_6t
Xbit_r102_c136 bl_136 br_136 wl_102 vdd gnd cell_6t
Xbit_r103_c136 bl_136 br_136 wl_103 vdd gnd cell_6t
Xbit_r104_c136 bl_136 br_136 wl_104 vdd gnd cell_6t
Xbit_r105_c136 bl_136 br_136 wl_105 vdd gnd cell_6t
Xbit_r106_c136 bl_136 br_136 wl_106 vdd gnd cell_6t
Xbit_r107_c136 bl_136 br_136 wl_107 vdd gnd cell_6t
Xbit_r108_c136 bl_136 br_136 wl_108 vdd gnd cell_6t
Xbit_r109_c136 bl_136 br_136 wl_109 vdd gnd cell_6t
Xbit_r110_c136 bl_136 br_136 wl_110 vdd gnd cell_6t
Xbit_r111_c136 bl_136 br_136 wl_111 vdd gnd cell_6t
Xbit_r112_c136 bl_136 br_136 wl_112 vdd gnd cell_6t
Xbit_r113_c136 bl_136 br_136 wl_113 vdd gnd cell_6t
Xbit_r114_c136 bl_136 br_136 wl_114 vdd gnd cell_6t
Xbit_r115_c136 bl_136 br_136 wl_115 vdd gnd cell_6t
Xbit_r116_c136 bl_136 br_136 wl_116 vdd gnd cell_6t
Xbit_r117_c136 bl_136 br_136 wl_117 vdd gnd cell_6t
Xbit_r118_c136 bl_136 br_136 wl_118 vdd gnd cell_6t
Xbit_r119_c136 bl_136 br_136 wl_119 vdd gnd cell_6t
Xbit_r120_c136 bl_136 br_136 wl_120 vdd gnd cell_6t
Xbit_r121_c136 bl_136 br_136 wl_121 vdd gnd cell_6t
Xbit_r122_c136 bl_136 br_136 wl_122 vdd gnd cell_6t
Xbit_r123_c136 bl_136 br_136 wl_123 vdd gnd cell_6t
Xbit_r124_c136 bl_136 br_136 wl_124 vdd gnd cell_6t
Xbit_r125_c136 bl_136 br_136 wl_125 vdd gnd cell_6t
Xbit_r126_c136 bl_136 br_136 wl_126 vdd gnd cell_6t
Xbit_r127_c136 bl_136 br_136 wl_127 vdd gnd cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd cell_6t
Xbit_r1_c137 bl_137 br_137 wl_1 vdd gnd cell_6t
Xbit_r2_c137 bl_137 br_137 wl_2 vdd gnd cell_6t
Xbit_r3_c137 bl_137 br_137 wl_3 vdd gnd cell_6t
Xbit_r4_c137 bl_137 br_137 wl_4 vdd gnd cell_6t
Xbit_r5_c137 bl_137 br_137 wl_5 vdd gnd cell_6t
Xbit_r6_c137 bl_137 br_137 wl_6 vdd gnd cell_6t
Xbit_r7_c137 bl_137 br_137 wl_7 vdd gnd cell_6t
Xbit_r8_c137 bl_137 br_137 wl_8 vdd gnd cell_6t
Xbit_r9_c137 bl_137 br_137 wl_9 vdd gnd cell_6t
Xbit_r10_c137 bl_137 br_137 wl_10 vdd gnd cell_6t
Xbit_r11_c137 bl_137 br_137 wl_11 vdd gnd cell_6t
Xbit_r12_c137 bl_137 br_137 wl_12 vdd gnd cell_6t
Xbit_r13_c137 bl_137 br_137 wl_13 vdd gnd cell_6t
Xbit_r14_c137 bl_137 br_137 wl_14 vdd gnd cell_6t
Xbit_r15_c137 bl_137 br_137 wl_15 vdd gnd cell_6t
Xbit_r16_c137 bl_137 br_137 wl_16 vdd gnd cell_6t
Xbit_r17_c137 bl_137 br_137 wl_17 vdd gnd cell_6t
Xbit_r18_c137 bl_137 br_137 wl_18 vdd gnd cell_6t
Xbit_r19_c137 bl_137 br_137 wl_19 vdd gnd cell_6t
Xbit_r20_c137 bl_137 br_137 wl_20 vdd gnd cell_6t
Xbit_r21_c137 bl_137 br_137 wl_21 vdd gnd cell_6t
Xbit_r22_c137 bl_137 br_137 wl_22 vdd gnd cell_6t
Xbit_r23_c137 bl_137 br_137 wl_23 vdd gnd cell_6t
Xbit_r24_c137 bl_137 br_137 wl_24 vdd gnd cell_6t
Xbit_r25_c137 bl_137 br_137 wl_25 vdd gnd cell_6t
Xbit_r26_c137 bl_137 br_137 wl_26 vdd gnd cell_6t
Xbit_r27_c137 bl_137 br_137 wl_27 vdd gnd cell_6t
Xbit_r28_c137 bl_137 br_137 wl_28 vdd gnd cell_6t
Xbit_r29_c137 bl_137 br_137 wl_29 vdd gnd cell_6t
Xbit_r30_c137 bl_137 br_137 wl_30 vdd gnd cell_6t
Xbit_r31_c137 bl_137 br_137 wl_31 vdd gnd cell_6t
Xbit_r32_c137 bl_137 br_137 wl_32 vdd gnd cell_6t
Xbit_r33_c137 bl_137 br_137 wl_33 vdd gnd cell_6t
Xbit_r34_c137 bl_137 br_137 wl_34 vdd gnd cell_6t
Xbit_r35_c137 bl_137 br_137 wl_35 vdd gnd cell_6t
Xbit_r36_c137 bl_137 br_137 wl_36 vdd gnd cell_6t
Xbit_r37_c137 bl_137 br_137 wl_37 vdd gnd cell_6t
Xbit_r38_c137 bl_137 br_137 wl_38 vdd gnd cell_6t
Xbit_r39_c137 bl_137 br_137 wl_39 vdd gnd cell_6t
Xbit_r40_c137 bl_137 br_137 wl_40 vdd gnd cell_6t
Xbit_r41_c137 bl_137 br_137 wl_41 vdd gnd cell_6t
Xbit_r42_c137 bl_137 br_137 wl_42 vdd gnd cell_6t
Xbit_r43_c137 bl_137 br_137 wl_43 vdd gnd cell_6t
Xbit_r44_c137 bl_137 br_137 wl_44 vdd gnd cell_6t
Xbit_r45_c137 bl_137 br_137 wl_45 vdd gnd cell_6t
Xbit_r46_c137 bl_137 br_137 wl_46 vdd gnd cell_6t
Xbit_r47_c137 bl_137 br_137 wl_47 vdd gnd cell_6t
Xbit_r48_c137 bl_137 br_137 wl_48 vdd gnd cell_6t
Xbit_r49_c137 bl_137 br_137 wl_49 vdd gnd cell_6t
Xbit_r50_c137 bl_137 br_137 wl_50 vdd gnd cell_6t
Xbit_r51_c137 bl_137 br_137 wl_51 vdd gnd cell_6t
Xbit_r52_c137 bl_137 br_137 wl_52 vdd gnd cell_6t
Xbit_r53_c137 bl_137 br_137 wl_53 vdd gnd cell_6t
Xbit_r54_c137 bl_137 br_137 wl_54 vdd gnd cell_6t
Xbit_r55_c137 bl_137 br_137 wl_55 vdd gnd cell_6t
Xbit_r56_c137 bl_137 br_137 wl_56 vdd gnd cell_6t
Xbit_r57_c137 bl_137 br_137 wl_57 vdd gnd cell_6t
Xbit_r58_c137 bl_137 br_137 wl_58 vdd gnd cell_6t
Xbit_r59_c137 bl_137 br_137 wl_59 vdd gnd cell_6t
Xbit_r60_c137 bl_137 br_137 wl_60 vdd gnd cell_6t
Xbit_r61_c137 bl_137 br_137 wl_61 vdd gnd cell_6t
Xbit_r62_c137 bl_137 br_137 wl_62 vdd gnd cell_6t
Xbit_r63_c137 bl_137 br_137 wl_63 vdd gnd cell_6t
Xbit_r64_c137 bl_137 br_137 wl_64 vdd gnd cell_6t
Xbit_r65_c137 bl_137 br_137 wl_65 vdd gnd cell_6t
Xbit_r66_c137 bl_137 br_137 wl_66 vdd gnd cell_6t
Xbit_r67_c137 bl_137 br_137 wl_67 vdd gnd cell_6t
Xbit_r68_c137 bl_137 br_137 wl_68 vdd gnd cell_6t
Xbit_r69_c137 bl_137 br_137 wl_69 vdd gnd cell_6t
Xbit_r70_c137 bl_137 br_137 wl_70 vdd gnd cell_6t
Xbit_r71_c137 bl_137 br_137 wl_71 vdd gnd cell_6t
Xbit_r72_c137 bl_137 br_137 wl_72 vdd gnd cell_6t
Xbit_r73_c137 bl_137 br_137 wl_73 vdd gnd cell_6t
Xbit_r74_c137 bl_137 br_137 wl_74 vdd gnd cell_6t
Xbit_r75_c137 bl_137 br_137 wl_75 vdd gnd cell_6t
Xbit_r76_c137 bl_137 br_137 wl_76 vdd gnd cell_6t
Xbit_r77_c137 bl_137 br_137 wl_77 vdd gnd cell_6t
Xbit_r78_c137 bl_137 br_137 wl_78 vdd gnd cell_6t
Xbit_r79_c137 bl_137 br_137 wl_79 vdd gnd cell_6t
Xbit_r80_c137 bl_137 br_137 wl_80 vdd gnd cell_6t
Xbit_r81_c137 bl_137 br_137 wl_81 vdd gnd cell_6t
Xbit_r82_c137 bl_137 br_137 wl_82 vdd gnd cell_6t
Xbit_r83_c137 bl_137 br_137 wl_83 vdd gnd cell_6t
Xbit_r84_c137 bl_137 br_137 wl_84 vdd gnd cell_6t
Xbit_r85_c137 bl_137 br_137 wl_85 vdd gnd cell_6t
Xbit_r86_c137 bl_137 br_137 wl_86 vdd gnd cell_6t
Xbit_r87_c137 bl_137 br_137 wl_87 vdd gnd cell_6t
Xbit_r88_c137 bl_137 br_137 wl_88 vdd gnd cell_6t
Xbit_r89_c137 bl_137 br_137 wl_89 vdd gnd cell_6t
Xbit_r90_c137 bl_137 br_137 wl_90 vdd gnd cell_6t
Xbit_r91_c137 bl_137 br_137 wl_91 vdd gnd cell_6t
Xbit_r92_c137 bl_137 br_137 wl_92 vdd gnd cell_6t
Xbit_r93_c137 bl_137 br_137 wl_93 vdd gnd cell_6t
Xbit_r94_c137 bl_137 br_137 wl_94 vdd gnd cell_6t
Xbit_r95_c137 bl_137 br_137 wl_95 vdd gnd cell_6t
Xbit_r96_c137 bl_137 br_137 wl_96 vdd gnd cell_6t
Xbit_r97_c137 bl_137 br_137 wl_97 vdd gnd cell_6t
Xbit_r98_c137 bl_137 br_137 wl_98 vdd gnd cell_6t
Xbit_r99_c137 bl_137 br_137 wl_99 vdd gnd cell_6t
Xbit_r100_c137 bl_137 br_137 wl_100 vdd gnd cell_6t
Xbit_r101_c137 bl_137 br_137 wl_101 vdd gnd cell_6t
Xbit_r102_c137 bl_137 br_137 wl_102 vdd gnd cell_6t
Xbit_r103_c137 bl_137 br_137 wl_103 vdd gnd cell_6t
Xbit_r104_c137 bl_137 br_137 wl_104 vdd gnd cell_6t
Xbit_r105_c137 bl_137 br_137 wl_105 vdd gnd cell_6t
Xbit_r106_c137 bl_137 br_137 wl_106 vdd gnd cell_6t
Xbit_r107_c137 bl_137 br_137 wl_107 vdd gnd cell_6t
Xbit_r108_c137 bl_137 br_137 wl_108 vdd gnd cell_6t
Xbit_r109_c137 bl_137 br_137 wl_109 vdd gnd cell_6t
Xbit_r110_c137 bl_137 br_137 wl_110 vdd gnd cell_6t
Xbit_r111_c137 bl_137 br_137 wl_111 vdd gnd cell_6t
Xbit_r112_c137 bl_137 br_137 wl_112 vdd gnd cell_6t
Xbit_r113_c137 bl_137 br_137 wl_113 vdd gnd cell_6t
Xbit_r114_c137 bl_137 br_137 wl_114 vdd gnd cell_6t
Xbit_r115_c137 bl_137 br_137 wl_115 vdd gnd cell_6t
Xbit_r116_c137 bl_137 br_137 wl_116 vdd gnd cell_6t
Xbit_r117_c137 bl_137 br_137 wl_117 vdd gnd cell_6t
Xbit_r118_c137 bl_137 br_137 wl_118 vdd gnd cell_6t
Xbit_r119_c137 bl_137 br_137 wl_119 vdd gnd cell_6t
Xbit_r120_c137 bl_137 br_137 wl_120 vdd gnd cell_6t
Xbit_r121_c137 bl_137 br_137 wl_121 vdd gnd cell_6t
Xbit_r122_c137 bl_137 br_137 wl_122 vdd gnd cell_6t
Xbit_r123_c137 bl_137 br_137 wl_123 vdd gnd cell_6t
Xbit_r124_c137 bl_137 br_137 wl_124 vdd gnd cell_6t
Xbit_r125_c137 bl_137 br_137 wl_125 vdd gnd cell_6t
Xbit_r126_c137 bl_137 br_137 wl_126 vdd gnd cell_6t
Xbit_r127_c137 bl_137 br_137 wl_127 vdd gnd cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd cell_6t
Xbit_r1_c138 bl_138 br_138 wl_1 vdd gnd cell_6t
Xbit_r2_c138 bl_138 br_138 wl_2 vdd gnd cell_6t
Xbit_r3_c138 bl_138 br_138 wl_3 vdd gnd cell_6t
Xbit_r4_c138 bl_138 br_138 wl_4 vdd gnd cell_6t
Xbit_r5_c138 bl_138 br_138 wl_5 vdd gnd cell_6t
Xbit_r6_c138 bl_138 br_138 wl_6 vdd gnd cell_6t
Xbit_r7_c138 bl_138 br_138 wl_7 vdd gnd cell_6t
Xbit_r8_c138 bl_138 br_138 wl_8 vdd gnd cell_6t
Xbit_r9_c138 bl_138 br_138 wl_9 vdd gnd cell_6t
Xbit_r10_c138 bl_138 br_138 wl_10 vdd gnd cell_6t
Xbit_r11_c138 bl_138 br_138 wl_11 vdd gnd cell_6t
Xbit_r12_c138 bl_138 br_138 wl_12 vdd gnd cell_6t
Xbit_r13_c138 bl_138 br_138 wl_13 vdd gnd cell_6t
Xbit_r14_c138 bl_138 br_138 wl_14 vdd gnd cell_6t
Xbit_r15_c138 bl_138 br_138 wl_15 vdd gnd cell_6t
Xbit_r16_c138 bl_138 br_138 wl_16 vdd gnd cell_6t
Xbit_r17_c138 bl_138 br_138 wl_17 vdd gnd cell_6t
Xbit_r18_c138 bl_138 br_138 wl_18 vdd gnd cell_6t
Xbit_r19_c138 bl_138 br_138 wl_19 vdd gnd cell_6t
Xbit_r20_c138 bl_138 br_138 wl_20 vdd gnd cell_6t
Xbit_r21_c138 bl_138 br_138 wl_21 vdd gnd cell_6t
Xbit_r22_c138 bl_138 br_138 wl_22 vdd gnd cell_6t
Xbit_r23_c138 bl_138 br_138 wl_23 vdd gnd cell_6t
Xbit_r24_c138 bl_138 br_138 wl_24 vdd gnd cell_6t
Xbit_r25_c138 bl_138 br_138 wl_25 vdd gnd cell_6t
Xbit_r26_c138 bl_138 br_138 wl_26 vdd gnd cell_6t
Xbit_r27_c138 bl_138 br_138 wl_27 vdd gnd cell_6t
Xbit_r28_c138 bl_138 br_138 wl_28 vdd gnd cell_6t
Xbit_r29_c138 bl_138 br_138 wl_29 vdd gnd cell_6t
Xbit_r30_c138 bl_138 br_138 wl_30 vdd gnd cell_6t
Xbit_r31_c138 bl_138 br_138 wl_31 vdd gnd cell_6t
Xbit_r32_c138 bl_138 br_138 wl_32 vdd gnd cell_6t
Xbit_r33_c138 bl_138 br_138 wl_33 vdd gnd cell_6t
Xbit_r34_c138 bl_138 br_138 wl_34 vdd gnd cell_6t
Xbit_r35_c138 bl_138 br_138 wl_35 vdd gnd cell_6t
Xbit_r36_c138 bl_138 br_138 wl_36 vdd gnd cell_6t
Xbit_r37_c138 bl_138 br_138 wl_37 vdd gnd cell_6t
Xbit_r38_c138 bl_138 br_138 wl_38 vdd gnd cell_6t
Xbit_r39_c138 bl_138 br_138 wl_39 vdd gnd cell_6t
Xbit_r40_c138 bl_138 br_138 wl_40 vdd gnd cell_6t
Xbit_r41_c138 bl_138 br_138 wl_41 vdd gnd cell_6t
Xbit_r42_c138 bl_138 br_138 wl_42 vdd gnd cell_6t
Xbit_r43_c138 bl_138 br_138 wl_43 vdd gnd cell_6t
Xbit_r44_c138 bl_138 br_138 wl_44 vdd gnd cell_6t
Xbit_r45_c138 bl_138 br_138 wl_45 vdd gnd cell_6t
Xbit_r46_c138 bl_138 br_138 wl_46 vdd gnd cell_6t
Xbit_r47_c138 bl_138 br_138 wl_47 vdd gnd cell_6t
Xbit_r48_c138 bl_138 br_138 wl_48 vdd gnd cell_6t
Xbit_r49_c138 bl_138 br_138 wl_49 vdd gnd cell_6t
Xbit_r50_c138 bl_138 br_138 wl_50 vdd gnd cell_6t
Xbit_r51_c138 bl_138 br_138 wl_51 vdd gnd cell_6t
Xbit_r52_c138 bl_138 br_138 wl_52 vdd gnd cell_6t
Xbit_r53_c138 bl_138 br_138 wl_53 vdd gnd cell_6t
Xbit_r54_c138 bl_138 br_138 wl_54 vdd gnd cell_6t
Xbit_r55_c138 bl_138 br_138 wl_55 vdd gnd cell_6t
Xbit_r56_c138 bl_138 br_138 wl_56 vdd gnd cell_6t
Xbit_r57_c138 bl_138 br_138 wl_57 vdd gnd cell_6t
Xbit_r58_c138 bl_138 br_138 wl_58 vdd gnd cell_6t
Xbit_r59_c138 bl_138 br_138 wl_59 vdd gnd cell_6t
Xbit_r60_c138 bl_138 br_138 wl_60 vdd gnd cell_6t
Xbit_r61_c138 bl_138 br_138 wl_61 vdd gnd cell_6t
Xbit_r62_c138 bl_138 br_138 wl_62 vdd gnd cell_6t
Xbit_r63_c138 bl_138 br_138 wl_63 vdd gnd cell_6t
Xbit_r64_c138 bl_138 br_138 wl_64 vdd gnd cell_6t
Xbit_r65_c138 bl_138 br_138 wl_65 vdd gnd cell_6t
Xbit_r66_c138 bl_138 br_138 wl_66 vdd gnd cell_6t
Xbit_r67_c138 bl_138 br_138 wl_67 vdd gnd cell_6t
Xbit_r68_c138 bl_138 br_138 wl_68 vdd gnd cell_6t
Xbit_r69_c138 bl_138 br_138 wl_69 vdd gnd cell_6t
Xbit_r70_c138 bl_138 br_138 wl_70 vdd gnd cell_6t
Xbit_r71_c138 bl_138 br_138 wl_71 vdd gnd cell_6t
Xbit_r72_c138 bl_138 br_138 wl_72 vdd gnd cell_6t
Xbit_r73_c138 bl_138 br_138 wl_73 vdd gnd cell_6t
Xbit_r74_c138 bl_138 br_138 wl_74 vdd gnd cell_6t
Xbit_r75_c138 bl_138 br_138 wl_75 vdd gnd cell_6t
Xbit_r76_c138 bl_138 br_138 wl_76 vdd gnd cell_6t
Xbit_r77_c138 bl_138 br_138 wl_77 vdd gnd cell_6t
Xbit_r78_c138 bl_138 br_138 wl_78 vdd gnd cell_6t
Xbit_r79_c138 bl_138 br_138 wl_79 vdd gnd cell_6t
Xbit_r80_c138 bl_138 br_138 wl_80 vdd gnd cell_6t
Xbit_r81_c138 bl_138 br_138 wl_81 vdd gnd cell_6t
Xbit_r82_c138 bl_138 br_138 wl_82 vdd gnd cell_6t
Xbit_r83_c138 bl_138 br_138 wl_83 vdd gnd cell_6t
Xbit_r84_c138 bl_138 br_138 wl_84 vdd gnd cell_6t
Xbit_r85_c138 bl_138 br_138 wl_85 vdd gnd cell_6t
Xbit_r86_c138 bl_138 br_138 wl_86 vdd gnd cell_6t
Xbit_r87_c138 bl_138 br_138 wl_87 vdd gnd cell_6t
Xbit_r88_c138 bl_138 br_138 wl_88 vdd gnd cell_6t
Xbit_r89_c138 bl_138 br_138 wl_89 vdd gnd cell_6t
Xbit_r90_c138 bl_138 br_138 wl_90 vdd gnd cell_6t
Xbit_r91_c138 bl_138 br_138 wl_91 vdd gnd cell_6t
Xbit_r92_c138 bl_138 br_138 wl_92 vdd gnd cell_6t
Xbit_r93_c138 bl_138 br_138 wl_93 vdd gnd cell_6t
Xbit_r94_c138 bl_138 br_138 wl_94 vdd gnd cell_6t
Xbit_r95_c138 bl_138 br_138 wl_95 vdd gnd cell_6t
Xbit_r96_c138 bl_138 br_138 wl_96 vdd gnd cell_6t
Xbit_r97_c138 bl_138 br_138 wl_97 vdd gnd cell_6t
Xbit_r98_c138 bl_138 br_138 wl_98 vdd gnd cell_6t
Xbit_r99_c138 bl_138 br_138 wl_99 vdd gnd cell_6t
Xbit_r100_c138 bl_138 br_138 wl_100 vdd gnd cell_6t
Xbit_r101_c138 bl_138 br_138 wl_101 vdd gnd cell_6t
Xbit_r102_c138 bl_138 br_138 wl_102 vdd gnd cell_6t
Xbit_r103_c138 bl_138 br_138 wl_103 vdd gnd cell_6t
Xbit_r104_c138 bl_138 br_138 wl_104 vdd gnd cell_6t
Xbit_r105_c138 bl_138 br_138 wl_105 vdd gnd cell_6t
Xbit_r106_c138 bl_138 br_138 wl_106 vdd gnd cell_6t
Xbit_r107_c138 bl_138 br_138 wl_107 vdd gnd cell_6t
Xbit_r108_c138 bl_138 br_138 wl_108 vdd gnd cell_6t
Xbit_r109_c138 bl_138 br_138 wl_109 vdd gnd cell_6t
Xbit_r110_c138 bl_138 br_138 wl_110 vdd gnd cell_6t
Xbit_r111_c138 bl_138 br_138 wl_111 vdd gnd cell_6t
Xbit_r112_c138 bl_138 br_138 wl_112 vdd gnd cell_6t
Xbit_r113_c138 bl_138 br_138 wl_113 vdd gnd cell_6t
Xbit_r114_c138 bl_138 br_138 wl_114 vdd gnd cell_6t
Xbit_r115_c138 bl_138 br_138 wl_115 vdd gnd cell_6t
Xbit_r116_c138 bl_138 br_138 wl_116 vdd gnd cell_6t
Xbit_r117_c138 bl_138 br_138 wl_117 vdd gnd cell_6t
Xbit_r118_c138 bl_138 br_138 wl_118 vdd gnd cell_6t
Xbit_r119_c138 bl_138 br_138 wl_119 vdd gnd cell_6t
Xbit_r120_c138 bl_138 br_138 wl_120 vdd gnd cell_6t
Xbit_r121_c138 bl_138 br_138 wl_121 vdd gnd cell_6t
Xbit_r122_c138 bl_138 br_138 wl_122 vdd gnd cell_6t
Xbit_r123_c138 bl_138 br_138 wl_123 vdd gnd cell_6t
Xbit_r124_c138 bl_138 br_138 wl_124 vdd gnd cell_6t
Xbit_r125_c138 bl_138 br_138 wl_125 vdd gnd cell_6t
Xbit_r126_c138 bl_138 br_138 wl_126 vdd gnd cell_6t
Xbit_r127_c138 bl_138 br_138 wl_127 vdd gnd cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd cell_6t
Xbit_r1_c139 bl_139 br_139 wl_1 vdd gnd cell_6t
Xbit_r2_c139 bl_139 br_139 wl_2 vdd gnd cell_6t
Xbit_r3_c139 bl_139 br_139 wl_3 vdd gnd cell_6t
Xbit_r4_c139 bl_139 br_139 wl_4 vdd gnd cell_6t
Xbit_r5_c139 bl_139 br_139 wl_5 vdd gnd cell_6t
Xbit_r6_c139 bl_139 br_139 wl_6 vdd gnd cell_6t
Xbit_r7_c139 bl_139 br_139 wl_7 vdd gnd cell_6t
Xbit_r8_c139 bl_139 br_139 wl_8 vdd gnd cell_6t
Xbit_r9_c139 bl_139 br_139 wl_9 vdd gnd cell_6t
Xbit_r10_c139 bl_139 br_139 wl_10 vdd gnd cell_6t
Xbit_r11_c139 bl_139 br_139 wl_11 vdd gnd cell_6t
Xbit_r12_c139 bl_139 br_139 wl_12 vdd gnd cell_6t
Xbit_r13_c139 bl_139 br_139 wl_13 vdd gnd cell_6t
Xbit_r14_c139 bl_139 br_139 wl_14 vdd gnd cell_6t
Xbit_r15_c139 bl_139 br_139 wl_15 vdd gnd cell_6t
Xbit_r16_c139 bl_139 br_139 wl_16 vdd gnd cell_6t
Xbit_r17_c139 bl_139 br_139 wl_17 vdd gnd cell_6t
Xbit_r18_c139 bl_139 br_139 wl_18 vdd gnd cell_6t
Xbit_r19_c139 bl_139 br_139 wl_19 vdd gnd cell_6t
Xbit_r20_c139 bl_139 br_139 wl_20 vdd gnd cell_6t
Xbit_r21_c139 bl_139 br_139 wl_21 vdd gnd cell_6t
Xbit_r22_c139 bl_139 br_139 wl_22 vdd gnd cell_6t
Xbit_r23_c139 bl_139 br_139 wl_23 vdd gnd cell_6t
Xbit_r24_c139 bl_139 br_139 wl_24 vdd gnd cell_6t
Xbit_r25_c139 bl_139 br_139 wl_25 vdd gnd cell_6t
Xbit_r26_c139 bl_139 br_139 wl_26 vdd gnd cell_6t
Xbit_r27_c139 bl_139 br_139 wl_27 vdd gnd cell_6t
Xbit_r28_c139 bl_139 br_139 wl_28 vdd gnd cell_6t
Xbit_r29_c139 bl_139 br_139 wl_29 vdd gnd cell_6t
Xbit_r30_c139 bl_139 br_139 wl_30 vdd gnd cell_6t
Xbit_r31_c139 bl_139 br_139 wl_31 vdd gnd cell_6t
Xbit_r32_c139 bl_139 br_139 wl_32 vdd gnd cell_6t
Xbit_r33_c139 bl_139 br_139 wl_33 vdd gnd cell_6t
Xbit_r34_c139 bl_139 br_139 wl_34 vdd gnd cell_6t
Xbit_r35_c139 bl_139 br_139 wl_35 vdd gnd cell_6t
Xbit_r36_c139 bl_139 br_139 wl_36 vdd gnd cell_6t
Xbit_r37_c139 bl_139 br_139 wl_37 vdd gnd cell_6t
Xbit_r38_c139 bl_139 br_139 wl_38 vdd gnd cell_6t
Xbit_r39_c139 bl_139 br_139 wl_39 vdd gnd cell_6t
Xbit_r40_c139 bl_139 br_139 wl_40 vdd gnd cell_6t
Xbit_r41_c139 bl_139 br_139 wl_41 vdd gnd cell_6t
Xbit_r42_c139 bl_139 br_139 wl_42 vdd gnd cell_6t
Xbit_r43_c139 bl_139 br_139 wl_43 vdd gnd cell_6t
Xbit_r44_c139 bl_139 br_139 wl_44 vdd gnd cell_6t
Xbit_r45_c139 bl_139 br_139 wl_45 vdd gnd cell_6t
Xbit_r46_c139 bl_139 br_139 wl_46 vdd gnd cell_6t
Xbit_r47_c139 bl_139 br_139 wl_47 vdd gnd cell_6t
Xbit_r48_c139 bl_139 br_139 wl_48 vdd gnd cell_6t
Xbit_r49_c139 bl_139 br_139 wl_49 vdd gnd cell_6t
Xbit_r50_c139 bl_139 br_139 wl_50 vdd gnd cell_6t
Xbit_r51_c139 bl_139 br_139 wl_51 vdd gnd cell_6t
Xbit_r52_c139 bl_139 br_139 wl_52 vdd gnd cell_6t
Xbit_r53_c139 bl_139 br_139 wl_53 vdd gnd cell_6t
Xbit_r54_c139 bl_139 br_139 wl_54 vdd gnd cell_6t
Xbit_r55_c139 bl_139 br_139 wl_55 vdd gnd cell_6t
Xbit_r56_c139 bl_139 br_139 wl_56 vdd gnd cell_6t
Xbit_r57_c139 bl_139 br_139 wl_57 vdd gnd cell_6t
Xbit_r58_c139 bl_139 br_139 wl_58 vdd gnd cell_6t
Xbit_r59_c139 bl_139 br_139 wl_59 vdd gnd cell_6t
Xbit_r60_c139 bl_139 br_139 wl_60 vdd gnd cell_6t
Xbit_r61_c139 bl_139 br_139 wl_61 vdd gnd cell_6t
Xbit_r62_c139 bl_139 br_139 wl_62 vdd gnd cell_6t
Xbit_r63_c139 bl_139 br_139 wl_63 vdd gnd cell_6t
Xbit_r64_c139 bl_139 br_139 wl_64 vdd gnd cell_6t
Xbit_r65_c139 bl_139 br_139 wl_65 vdd gnd cell_6t
Xbit_r66_c139 bl_139 br_139 wl_66 vdd gnd cell_6t
Xbit_r67_c139 bl_139 br_139 wl_67 vdd gnd cell_6t
Xbit_r68_c139 bl_139 br_139 wl_68 vdd gnd cell_6t
Xbit_r69_c139 bl_139 br_139 wl_69 vdd gnd cell_6t
Xbit_r70_c139 bl_139 br_139 wl_70 vdd gnd cell_6t
Xbit_r71_c139 bl_139 br_139 wl_71 vdd gnd cell_6t
Xbit_r72_c139 bl_139 br_139 wl_72 vdd gnd cell_6t
Xbit_r73_c139 bl_139 br_139 wl_73 vdd gnd cell_6t
Xbit_r74_c139 bl_139 br_139 wl_74 vdd gnd cell_6t
Xbit_r75_c139 bl_139 br_139 wl_75 vdd gnd cell_6t
Xbit_r76_c139 bl_139 br_139 wl_76 vdd gnd cell_6t
Xbit_r77_c139 bl_139 br_139 wl_77 vdd gnd cell_6t
Xbit_r78_c139 bl_139 br_139 wl_78 vdd gnd cell_6t
Xbit_r79_c139 bl_139 br_139 wl_79 vdd gnd cell_6t
Xbit_r80_c139 bl_139 br_139 wl_80 vdd gnd cell_6t
Xbit_r81_c139 bl_139 br_139 wl_81 vdd gnd cell_6t
Xbit_r82_c139 bl_139 br_139 wl_82 vdd gnd cell_6t
Xbit_r83_c139 bl_139 br_139 wl_83 vdd gnd cell_6t
Xbit_r84_c139 bl_139 br_139 wl_84 vdd gnd cell_6t
Xbit_r85_c139 bl_139 br_139 wl_85 vdd gnd cell_6t
Xbit_r86_c139 bl_139 br_139 wl_86 vdd gnd cell_6t
Xbit_r87_c139 bl_139 br_139 wl_87 vdd gnd cell_6t
Xbit_r88_c139 bl_139 br_139 wl_88 vdd gnd cell_6t
Xbit_r89_c139 bl_139 br_139 wl_89 vdd gnd cell_6t
Xbit_r90_c139 bl_139 br_139 wl_90 vdd gnd cell_6t
Xbit_r91_c139 bl_139 br_139 wl_91 vdd gnd cell_6t
Xbit_r92_c139 bl_139 br_139 wl_92 vdd gnd cell_6t
Xbit_r93_c139 bl_139 br_139 wl_93 vdd gnd cell_6t
Xbit_r94_c139 bl_139 br_139 wl_94 vdd gnd cell_6t
Xbit_r95_c139 bl_139 br_139 wl_95 vdd gnd cell_6t
Xbit_r96_c139 bl_139 br_139 wl_96 vdd gnd cell_6t
Xbit_r97_c139 bl_139 br_139 wl_97 vdd gnd cell_6t
Xbit_r98_c139 bl_139 br_139 wl_98 vdd gnd cell_6t
Xbit_r99_c139 bl_139 br_139 wl_99 vdd gnd cell_6t
Xbit_r100_c139 bl_139 br_139 wl_100 vdd gnd cell_6t
Xbit_r101_c139 bl_139 br_139 wl_101 vdd gnd cell_6t
Xbit_r102_c139 bl_139 br_139 wl_102 vdd gnd cell_6t
Xbit_r103_c139 bl_139 br_139 wl_103 vdd gnd cell_6t
Xbit_r104_c139 bl_139 br_139 wl_104 vdd gnd cell_6t
Xbit_r105_c139 bl_139 br_139 wl_105 vdd gnd cell_6t
Xbit_r106_c139 bl_139 br_139 wl_106 vdd gnd cell_6t
Xbit_r107_c139 bl_139 br_139 wl_107 vdd gnd cell_6t
Xbit_r108_c139 bl_139 br_139 wl_108 vdd gnd cell_6t
Xbit_r109_c139 bl_139 br_139 wl_109 vdd gnd cell_6t
Xbit_r110_c139 bl_139 br_139 wl_110 vdd gnd cell_6t
Xbit_r111_c139 bl_139 br_139 wl_111 vdd gnd cell_6t
Xbit_r112_c139 bl_139 br_139 wl_112 vdd gnd cell_6t
Xbit_r113_c139 bl_139 br_139 wl_113 vdd gnd cell_6t
Xbit_r114_c139 bl_139 br_139 wl_114 vdd gnd cell_6t
Xbit_r115_c139 bl_139 br_139 wl_115 vdd gnd cell_6t
Xbit_r116_c139 bl_139 br_139 wl_116 vdd gnd cell_6t
Xbit_r117_c139 bl_139 br_139 wl_117 vdd gnd cell_6t
Xbit_r118_c139 bl_139 br_139 wl_118 vdd gnd cell_6t
Xbit_r119_c139 bl_139 br_139 wl_119 vdd gnd cell_6t
Xbit_r120_c139 bl_139 br_139 wl_120 vdd gnd cell_6t
Xbit_r121_c139 bl_139 br_139 wl_121 vdd gnd cell_6t
Xbit_r122_c139 bl_139 br_139 wl_122 vdd gnd cell_6t
Xbit_r123_c139 bl_139 br_139 wl_123 vdd gnd cell_6t
Xbit_r124_c139 bl_139 br_139 wl_124 vdd gnd cell_6t
Xbit_r125_c139 bl_139 br_139 wl_125 vdd gnd cell_6t
Xbit_r126_c139 bl_139 br_139 wl_126 vdd gnd cell_6t
Xbit_r127_c139 bl_139 br_139 wl_127 vdd gnd cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd cell_6t
Xbit_r1_c140 bl_140 br_140 wl_1 vdd gnd cell_6t
Xbit_r2_c140 bl_140 br_140 wl_2 vdd gnd cell_6t
Xbit_r3_c140 bl_140 br_140 wl_3 vdd gnd cell_6t
Xbit_r4_c140 bl_140 br_140 wl_4 vdd gnd cell_6t
Xbit_r5_c140 bl_140 br_140 wl_5 vdd gnd cell_6t
Xbit_r6_c140 bl_140 br_140 wl_6 vdd gnd cell_6t
Xbit_r7_c140 bl_140 br_140 wl_7 vdd gnd cell_6t
Xbit_r8_c140 bl_140 br_140 wl_8 vdd gnd cell_6t
Xbit_r9_c140 bl_140 br_140 wl_9 vdd gnd cell_6t
Xbit_r10_c140 bl_140 br_140 wl_10 vdd gnd cell_6t
Xbit_r11_c140 bl_140 br_140 wl_11 vdd gnd cell_6t
Xbit_r12_c140 bl_140 br_140 wl_12 vdd gnd cell_6t
Xbit_r13_c140 bl_140 br_140 wl_13 vdd gnd cell_6t
Xbit_r14_c140 bl_140 br_140 wl_14 vdd gnd cell_6t
Xbit_r15_c140 bl_140 br_140 wl_15 vdd gnd cell_6t
Xbit_r16_c140 bl_140 br_140 wl_16 vdd gnd cell_6t
Xbit_r17_c140 bl_140 br_140 wl_17 vdd gnd cell_6t
Xbit_r18_c140 bl_140 br_140 wl_18 vdd gnd cell_6t
Xbit_r19_c140 bl_140 br_140 wl_19 vdd gnd cell_6t
Xbit_r20_c140 bl_140 br_140 wl_20 vdd gnd cell_6t
Xbit_r21_c140 bl_140 br_140 wl_21 vdd gnd cell_6t
Xbit_r22_c140 bl_140 br_140 wl_22 vdd gnd cell_6t
Xbit_r23_c140 bl_140 br_140 wl_23 vdd gnd cell_6t
Xbit_r24_c140 bl_140 br_140 wl_24 vdd gnd cell_6t
Xbit_r25_c140 bl_140 br_140 wl_25 vdd gnd cell_6t
Xbit_r26_c140 bl_140 br_140 wl_26 vdd gnd cell_6t
Xbit_r27_c140 bl_140 br_140 wl_27 vdd gnd cell_6t
Xbit_r28_c140 bl_140 br_140 wl_28 vdd gnd cell_6t
Xbit_r29_c140 bl_140 br_140 wl_29 vdd gnd cell_6t
Xbit_r30_c140 bl_140 br_140 wl_30 vdd gnd cell_6t
Xbit_r31_c140 bl_140 br_140 wl_31 vdd gnd cell_6t
Xbit_r32_c140 bl_140 br_140 wl_32 vdd gnd cell_6t
Xbit_r33_c140 bl_140 br_140 wl_33 vdd gnd cell_6t
Xbit_r34_c140 bl_140 br_140 wl_34 vdd gnd cell_6t
Xbit_r35_c140 bl_140 br_140 wl_35 vdd gnd cell_6t
Xbit_r36_c140 bl_140 br_140 wl_36 vdd gnd cell_6t
Xbit_r37_c140 bl_140 br_140 wl_37 vdd gnd cell_6t
Xbit_r38_c140 bl_140 br_140 wl_38 vdd gnd cell_6t
Xbit_r39_c140 bl_140 br_140 wl_39 vdd gnd cell_6t
Xbit_r40_c140 bl_140 br_140 wl_40 vdd gnd cell_6t
Xbit_r41_c140 bl_140 br_140 wl_41 vdd gnd cell_6t
Xbit_r42_c140 bl_140 br_140 wl_42 vdd gnd cell_6t
Xbit_r43_c140 bl_140 br_140 wl_43 vdd gnd cell_6t
Xbit_r44_c140 bl_140 br_140 wl_44 vdd gnd cell_6t
Xbit_r45_c140 bl_140 br_140 wl_45 vdd gnd cell_6t
Xbit_r46_c140 bl_140 br_140 wl_46 vdd gnd cell_6t
Xbit_r47_c140 bl_140 br_140 wl_47 vdd gnd cell_6t
Xbit_r48_c140 bl_140 br_140 wl_48 vdd gnd cell_6t
Xbit_r49_c140 bl_140 br_140 wl_49 vdd gnd cell_6t
Xbit_r50_c140 bl_140 br_140 wl_50 vdd gnd cell_6t
Xbit_r51_c140 bl_140 br_140 wl_51 vdd gnd cell_6t
Xbit_r52_c140 bl_140 br_140 wl_52 vdd gnd cell_6t
Xbit_r53_c140 bl_140 br_140 wl_53 vdd gnd cell_6t
Xbit_r54_c140 bl_140 br_140 wl_54 vdd gnd cell_6t
Xbit_r55_c140 bl_140 br_140 wl_55 vdd gnd cell_6t
Xbit_r56_c140 bl_140 br_140 wl_56 vdd gnd cell_6t
Xbit_r57_c140 bl_140 br_140 wl_57 vdd gnd cell_6t
Xbit_r58_c140 bl_140 br_140 wl_58 vdd gnd cell_6t
Xbit_r59_c140 bl_140 br_140 wl_59 vdd gnd cell_6t
Xbit_r60_c140 bl_140 br_140 wl_60 vdd gnd cell_6t
Xbit_r61_c140 bl_140 br_140 wl_61 vdd gnd cell_6t
Xbit_r62_c140 bl_140 br_140 wl_62 vdd gnd cell_6t
Xbit_r63_c140 bl_140 br_140 wl_63 vdd gnd cell_6t
Xbit_r64_c140 bl_140 br_140 wl_64 vdd gnd cell_6t
Xbit_r65_c140 bl_140 br_140 wl_65 vdd gnd cell_6t
Xbit_r66_c140 bl_140 br_140 wl_66 vdd gnd cell_6t
Xbit_r67_c140 bl_140 br_140 wl_67 vdd gnd cell_6t
Xbit_r68_c140 bl_140 br_140 wl_68 vdd gnd cell_6t
Xbit_r69_c140 bl_140 br_140 wl_69 vdd gnd cell_6t
Xbit_r70_c140 bl_140 br_140 wl_70 vdd gnd cell_6t
Xbit_r71_c140 bl_140 br_140 wl_71 vdd gnd cell_6t
Xbit_r72_c140 bl_140 br_140 wl_72 vdd gnd cell_6t
Xbit_r73_c140 bl_140 br_140 wl_73 vdd gnd cell_6t
Xbit_r74_c140 bl_140 br_140 wl_74 vdd gnd cell_6t
Xbit_r75_c140 bl_140 br_140 wl_75 vdd gnd cell_6t
Xbit_r76_c140 bl_140 br_140 wl_76 vdd gnd cell_6t
Xbit_r77_c140 bl_140 br_140 wl_77 vdd gnd cell_6t
Xbit_r78_c140 bl_140 br_140 wl_78 vdd gnd cell_6t
Xbit_r79_c140 bl_140 br_140 wl_79 vdd gnd cell_6t
Xbit_r80_c140 bl_140 br_140 wl_80 vdd gnd cell_6t
Xbit_r81_c140 bl_140 br_140 wl_81 vdd gnd cell_6t
Xbit_r82_c140 bl_140 br_140 wl_82 vdd gnd cell_6t
Xbit_r83_c140 bl_140 br_140 wl_83 vdd gnd cell_6t
Xbit_r84_c140 bl_140 br_140 wl_84 vdd gnd cell_6t
Xbit_r85_c140 bl_140 br_140 wl_85 vdd gnd cell_6t
Xbit_r86_c140 bl_140 br_140 wl_86 vdd gnd cell_6t
Xbit_r87_c140 bl_140 br_140 wl_87 vdd gnd cell_6t
Xbit_r88_c140 bl_140 br_140 wl_88 vdd gnd cell_6t
Xbit_r89_c140 bl_140 br_140 wl_89 vdd gnd cell_6t
Xbit_r90_c140 bl_140 br_140 wl_90 vdd gnd cell_6t
Xbit_r91_c140 bl_140 br_140 wl_91 vdd gnd cell_6t
Xbit_r92_c140 bl_140 br_140 wl_92 vdd gnd cell_6t
Xbit_r93_c140 bl_140 br_140 wl_93 vdd gnd cell_6t
Xbit_r94_c140 bl_140 br_140 wl_94 vdd gnd cell_6t
Xbit_r95_c140 bl_140 br_140 wl_95 vdd gnd cell_6t
Xbit_r96_c140 bl_140 br_140 wl_96 vdd gnd cell_6t
Xbit_r97_c140 bl_140 br_140 wl_97 vdd gnd cell_6t
Xbit_r98_c140 bl_140 br_140 wl_98 vdd gnd cell_6t
Xbit_r99_c140 bl_140 br_140 wl_99 vdd gnd cell_6t
Xbit_r100_c140 bl_140 br_140 wl_100 vdd gnd cell_6t
Xbit_r101_c140 bl_140 br_140 wl_101 vdd gnd cell_6t
Xbit_r102_c140 bl_140 br_140 wl_102 vdd gnd cell_6t
Xbit_r103_c140 bl_140 br_140 wl_103 vdd gnd cell_6t
Xbit_r104_c140 bl_140 br_140 wl_104 vdd gnd cell_6t
Xbit_r105_c140 bl_140 br_140 wl_105 vdd gnd cell_6t
Xbit_r106_c140 bl_140 br_140 wl_106 vdd gnd cell_6t
Xbit_r107_c140 bl_140 br_140 wl_107 vdd gnd cell_6t
Xbit_r108_c140 bl_140 br_140 wl_108 vdd gnd cell_6t
Xbit_r109_c140 bl_140 br_140 wl_109 vdd gnd cell_6t
Xbit_r110_c140 bl_140 br_140 wl_110 vdd gnd cell_6t
Xbit_r111_c140 bl_140 br_140 wl_111 vdd gnd cell_6t
Xbit_r112_c140 bl_140 br_140 wl_112 vdd gnd cell_6t
Xbit_r113_c140 bl_140 br_140 wl_113 vdd gnd cell_6t
Xbit_r114_c140 bl_140 br_140 wl_114 vdd gnd cell_6t
Xbit_r115_c140 bl_140 br_140 wl_115 vdd gnd cell_6t
Xbit_r116_c140 bl_140 br_140 wl_116 vdd gnd cell_6t
Xbit_r117_c140 bl_140 br_140 wl_117 vdd gnd cell_6t
Xbit_r118_c140 bl_140 br_140 wl_118 vdd gnd cell_6t
Xbit_r119_c140 bl_140 br_140 wl_119 vdd gnd cell_6t
Xbit_r120_c140 bl_140 br_140 wl_120 vdd gnd cell_6t
Xbit_r121_c140 bl_140 br_140 wl_121 vdd gnd cell_6t
Xbit_r122_c140 bl_140 br_140 wl_122 vdd gnd cell_6t
Xbit_r123_c140 bl_140 br_140 wl_123 vdd gnd cell_6t
Xbit_r124_c140 bl_140 br_140 wl_124 vdd gnd cell_6t
Xbit_r125_c140 bl_140 br_140 wl_125 vdd gnd cell_6t
Xbit_r126_c140 bl_140 br_140 wl_126 vdd gnd cell_6t
Xbit_r127_c140 bl_140 br_140 wl_127 vdd gnd cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd cell_6t
Xbit_r1_c141 bl_141 br_141 wl_1 vdd gnd cell_6t
Xbit_r2_c141 bl_141 br_141 wl_2 vdd gnd cell_6t
Xbit_r3_c141 bl_141 br_141 wl_3 vdd gnd cell_6t
Xbit_r4_c141 bl_141 br_141 wl_4 vdd gnd cell_6t
Xbit_r5_c141 bl_141 br_141 wl_5 vdd gnd cell_6t
Xbit_r6_c141 bl_141 br_141 wl_6 vdd gnd cell_6t
Xbit_r7_c141 bl_141 br_141 wl_7 vdd gnd cell_6t
Xbit_r8_c141 bl_141 br_141 wl_8 vdd gnd cell_6t
Xbit_r9_c141 bl_141 br_141 wl_9 vdd gnd cell_6t
Xbit_r10_c141 bl_141 br_141 wl_10 vdd gnd cell_6t
Xbit_r11_c141 bl_141 br_141 wl_11 vdd gnd cell_6t
Xbit_r12_c141 bl_141 br_141 wl_12 vdd gnd cell_6t
Xbit_r13_c141 bl_141 br_141 wl_13 vdd gnd cell_6t
Xbit_r14_c141 bl_141 br_141 wl_14 vdd gnd cell_6t
Xbit_r15_c141 bl_141 br_141 wl_15 vdd gnd cell_6t
Xbit_r16_c141 bl_141 br_141 wl_16 vdd gnd cell_6t
Xbit_r17_c141 bl_141 br_141 wl_17 vdd gnd cell_6t
Xbit_r18_c141 bl_141 br_141 wl_18 vdd gnd cell_6t
Xbit_r19_c141 bl_141 br_141 wl_19 vdd gnd cell_6t
Xbit_r20_c141 bl_141 br_141 wl_20 vdd gnd cell_6t
Xbit_r21_c141 bl_141 br_141 wl_21 vdd gnd cell_6t
Xbit_r22_c141 bl_141 br_141 wl_22 vdd gnd cell_6t
Xbit_r23_c141 bl_141 br_141 wl_23 vdd gnd cell_6t
Xbit_r24_c141 bl_141 br_141 wl_24 vdd gnd cell_6t
Xbit_r25_c141 bl_141 br_141 wl_25 vdd gnd cell_6t
Xbit_r26_c141 bl_141 br_141 wl_26 vdd gnd cell_6t
Xbit_r27_c141 bl_141 br_141 wl_27 vdd gnd cell_6t
Xbit_r28_c141 bl_141 br_141 wl_28 vdd gnd cell_6t
Xbit_r29_c141 bl_141 br_141 wl_29 vdd gnd cell_6t
Xbit_r30_c141 bl_141 br_141 wl_30 vdd gnd cell_6t
Xbit_r31_c141 bl_141 br_141 wl_31 vdd gnd cell_6t
Xbit_r32_c141 bl_141 br_141 wl_32 vdd gnd cell_6t
Xbit_r33_c141 bl_141 br_141 wl_33 vdd gnd cell_6t
Xbit_r34_c141 bl_141 br_141 wl_34 vdd gnd cell_6t
Xbit_r35_c141 bl_141 br_141 wl_35 vdd gnd cell_6t
Xbit_r36_c141 bl_141 br_141 wl_36 vdd gnd cell_6t
Xbit_r37_c141 bl_141 br_141 wl_37 vdd gnd cell_6t
Xbit_r38_c141 bl_141 br_141 wl_38 vdd gnd cell_6t
Xbit_r39_c141 bl_141 br_141 wl_39 vdd gnd cell_6t
Xbit_r40_c141 bl_141 br_141 wl_40 vdd gnd cell_6t
Xbit_r41_c141 bl_141 br_141 wl_41 vdd gnd cell_6t
Xbit_r42_c141 bl_141 br_141 wl_42 vdd gnd cell_6t
Xbit_r43_c141 bl_141 br_141 wl_43 vdd gnd cell_6t
Xbit_r44_c141 bl_141 br_141 wl_44 vdd gnd cell_6t
Xbit_r45_c141 bl_141 br_141 wl_45 vdd gnd cell_6t
Xbit_r46_c141 bl_141 br_141 wl_46 vdd gnd cell_6t
Xbit_r47_c141 bl_141 br_141 wl_47 vdd gnd cell_6t
Xbit_r48_c141 bl_141 br_141 wl_48 vdd gnd cell_6t
Xbit_r49_c141 bl_141 br_141 wl_49 vdd gnd cell_6t
Xbit_r50_c141 bl_141 br_141 wl_50 vdd gnd cell_6t
Xbit_r51_c141 bl_141 br_141 wl_51 vdd gnd cell_6t
Xbit_r52_c141 bl_141 br_141 wl_52 vdd gnd cell_6t
Xbit_r53_c141 bl_141 br_141 wl_53 vdd gnd cell_6t
Xbit_r54_c141 bl_141 br_141 wl_54 vdd gnd cell_6t
Xbit_r55_c141 bl_141 br_141 wl_55 vdd gnd cell_6t
Xbit_r56_c141 bl_141 br_141 wl_56 vdd gnd cell_6t
Xbit_r57_c141 bl_141 br_141 wl_57 vdd gnd cell_6t
Xbit_r58_c141 bl_141 br_141 wl_58 vdd gnd cell_6t
Xbit_r59_c141 bl_141 br_141 wl_59 vdd gnd cell_6t
Xbit_r60_c141 bl_141 br_141 wl_60 vdd gnd cell_6t
Xbit_r61_c141 bl_141 br_141 wl_61 vdd gnd cell_6t
Xbit_r62_c141 bl_141 br_141 wl_62 vdd gnd cell_6t
Xbit_r63_c141 bl_141 br_141 wl_63 vdd gnd cell_6t
Xbit_r64_c141 bl_141 br_141 wl_64 vdd gnd cell_6t
Xbit_r65_c141 bl_141 br_141 wl_65 vdd gnd cell_6t
Xbit_r66_c141 bl_141 br_141 wl_66 vdd gnd cell_6t
Xbit_r67_c141 bl_141 br_141 wl_67 vdd gnd cell_6t
Xbit_r68_c141 bl_141 br_141 wl_68 vdd gnd cell_6t
Xbit_r69_c141 bl_141 br_141 wl_69 vdd gnd cell_6t
Xbit_r70_c141 bl_141 br_141 wl_70 vdd gnd cell_6t
Xbit_r71_c141 bl_141 br_141 wl_71 vdd gnd cell_6t
Xbit_r72_c141 bl_141 br_141 wl_72 vdd gnd cell_6t
Xbit_r73_c141 bl_141 br_141 wl_73 vdd gnd cell_6t
Xbit_r74_c141 bl_141 br_141 wl_74 vdd gnd cell_6t
Xbit_r75_c141 bl_141 br_141 wl_75 vdd gnd cell_6t
Xbit_r76_c141 bl_141 br_141 wl_76 vdd gnd cell_6t
Xbit_r77_c141 bl_141 br_141 wl_77 vdd gnd cell_6t
Xbit_r78_c141 bl_141 br_141 wl_78 vdd gnd cell_6t
Xbit_r79_c141 bl_141 br_141 wl_79 vdd gnd cell_6t
Xbit_r80_c141 bl_141 br_141 wl_80 vdd gnd cell_6t
Xbit_r81_c141 bl_141 br_141 wl_81 vdd gnd cell_6t
Xbit_r82_c141 bl_141 br_141 wl_82 vdd gnd cell_6t
Xbit_r83_c141 bl_141 br_141 wl_83 vdd gnd cell_6t
Xbit_r84_c141 bl_141 br_141 wl_84 vdd gnd cell_6t
Xbit_r85_c141 bl_141 br_141 wl_85 vdd gnd cell_6t
Xbit_r86_c141 bl_141 br_141 wl_86 vdd gnd cell_6t
Xbit_r87_c141 bl_141 br_141 wl_87 vdd gnd cell_6t
Xbit_r88_c141 bl_141 br_141 wl_88 vdd gnd cell_6t
Xbit_r89_c141 bl_141 br_141 wl_89 vdd gnd cell_6t
Xbit_r90_c141 bl_141 br_141 wl_90 vdd gnd cell_6t
Xbit_r91_c141 bl_141 br_141 wl_91 vdd gnd cell_6t
Xbit_r92_c141 bl_141 br_141 wl_92 vdd gnd cell_6t
Xbit_r93_c141 bl_141 br_141 wl_93 vdd gnd cell_6t
Xbit_r94_c141 bl_141 br_141 wl_94 vdd gnd cell_6t
Xbit_r95_c141 bl_141 br_141 wl_95 vdd gnd cell_6t
Xbit_r96_c141 bl_141 br_141 wl_96 vdd gnd cell_6t
Xbit_r97_c141 bl_141 br_141 wl_97 vdd gnd cell_6t
Xbit_r98_c141 bl_141 br_141 wl_98 vdd gnd cell_6t
Xbit_r99_c141 bl_141 br_141 wl_99 vdd gnd cell_6t
Xbit_r100_c141 bl_141 br_141 wl_100 vdd gnd cell_6t
Xbit_r101_c141 bl_141 br_141 wl_101 vdd gnd cell_6t
Xbit_r102_c141 bl_141 br_141 wl_102 vdd gnd cell_6t
Xbit_r103_c141 bl_141 br_141 wl_103 vdd gnd cell_6t
Xbit_r104_c141 bl_141 br_141 wl_104 vdd gnd cell_6t
Xbit_r105_c141 bl_141 br_141 wl_105 vdd gnd cell_6t
Xbit_r106_c141 bl_141 br_141 wl_106 vdd gnd cell_6t
Xbit_r107_c141 bl_141 br_141 wl_107 vdd gnd cell_6t
Xbit_r108_c141 bl_141 br_141 wl_108 vdd gnd cell_6t
Xbit_r109_c141 bl_141 br_141 wl_109 vdd gnd cell_6t
Xbit_r110_c141 bl_141 br_141 wl_110 vdd gnd cell_6t
Xbit_r111_c141 bl_141 br_141 wl_111 vdd gnd cell_6t
Xbit_r112_c141 bl_141 br_141 wl_112 vdd gnd cell_6t
Xbit_r113_c141 bl_141 br_141 wl_113 vdd gnd cell_6t
Xbit_r114_c141 bl_141 br_141 wl_114 vdd gnd cell_6t
Xbit_r115_c141 bl_141 br_141 wl_115 vdd gnd cell_6t
Xbit_r116_c141 bl_141 br_141 wl_116 vdd gnd cell_6t
Xbit_r117_c141 bl_141 br_141 wl_117 vdd gnd cell_6t
Xbit_r118_c141 bl_141 br_141 wl_118 vdd gnd cell_6t
Xbit_r119_c141 bl_141 br_141 wl_119 vdd gnd cell_6t
Xbit_r120_c141 bl_141 br_141 wl_120 vdd gnd cell_6t
Xbit_r121_c141 bl_141 br_141 wl_121 vdd gnd cell_6t
Xbit_r122_c141 bl_141 br_141 wl_122 vdd gnd cell_6t
Xbit_r123_c141 bl_141 br_141 wl_123 vdd gnd cell_6t
Xbit_r124_c141 bl_141 br_141 wl_124 vdd gnd cell_6t
Xbit_r125_c141 bl_141 br_141 wl_125 vdd gnd cell_6t
Xbit_r126_c141 bl_141 br_141 wl_126 vdd gnd cell_6t
Xbit_r127_c141 bl_141 br_141 wl_127 vdd gnd cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd cell_6t
Xbit_r1_c142 bl_142 br_142 wl_1 vdd gnd cell_6t
Xbit_r2_c142 bl_142 br_142 wl_2 vdd gnd cell_6t
Xbit_r3_c142 bl_142 br_142 wl_3 vdd gnd cell_6t
Xbit_r4_c142 bl_142 br_142 wl_4 vdd gnd cell_6t
Xbit_r5_c142 bl_142 br_142 wl_5 vdd gnd cell_6t
Xbit_r6_c142 bl_142 br_142 wl_6 vdd gnd cell_6t
Xbit_r7_c142 bl_142 br_142 wl_7 vdd gnd cell_6t
Xbit_r8_c142 bl_142 br_142 wl_8 vdd gnd cell_6t
Xbit_r9_c142 bl_142 br_142 wl_9 vdd gnd cell_6t
Xbit_r10_c142 bl_142 br_142 wl_10 vdd gnd cell_6t
Xbit_r11_c142 bl_142 br_142 wl_11 vdd gnd cell_6t
Xbit_r12_c142 bl_142 br_142 wl_12 vdd gnd cell_6t
Xbit_r13_c142 bl_142 br_142 wl_13 vdd gnd cell_6t
Xbit_r14_c142 bl_142 br_142 wl_14 vdd gnd cell_6t
Xbit_r15_c142 bl_142 br_142 wl_15 vdd gnd cell_6t
Xbit_r16_c142 bl_142 br_142 wl_16 vdd gnd cell_6t
Xbit_r17_c142 bl_142 br_142 wl_17 vdd gnd cell_6t
Xbit_r18_c142 bl_142 br_142 wl_18 vdd gnd cell_6t
Xbit_r19_c142 bl_142 br_142 wl_19 vdd gnd cell_6t
Xbit_r20_c142 bl_142 br_142 wl_20 vdd gnd cell_6t
Xbit_r21_c142 bl_142 br_142 wl_21 vdd gnd cell_6t
Xbit_r22_c142 bl_142 br_142 wl_22 vdd gnd cell_6t
Xbit_r23_c142 bl_142 br_142 wl_23 vdd gnd cell_6t
Xbit_r24_c142 bl_142 br_142 wl_24 vdd gnd cell_6t
Xbit_r25_c142 bl_142 br_142 wl_25 vdd gnd cell_6t
Xbit_r26_c142 bl_142 br_142 wl_26 vdd gnd cell_6t
Xbit_r27_c142 bl_142 br_142 wl_27 vdd gnd cell_6t
Xbit_r28_c142 bl_142 br_142 wl_28 vdd gnd cell_6t
Xbit_r29_c142 bl_142 br_142 wl_29 vdd gnd cell_6t
Xbit_r30_c142 bl_142 br_142 wl_30 vdd gnd cell_6t
Xbit_r31_c142 bl_142 br_142 wl_31 vdd gnd cell_6t
Xbit_r32_c142 bl_142 br_142 wl_32 vdd gnd cell_6t
Xbit_r33_c142 bl_142 br_142 wl_33 vdd gnd cell_6t
Xbit_r34_c142 bl_142 br_142 wl_34 vdd gnd cell_6t
Xbit_r35_c142 bl_142 br_142 wl_35 vdd gnd cell_6t
Xbit_r36_c142 bl_142 br_142 wl_36 vdd gnd cell_6t
Xbit_r37_c142 bl_142 br_142 wl_37 vdd gnd cell_6t
Xbit_r38_c142 bl_142 br_142 wl_38 vdd gnd cell_6t
Xbit_r39_c142 bl_142 br_142 wl_39 vdd gnd cell_6t
Xbit_r40_c142 bl_142 br_142 wl_40 vdd gnd cell_6t
Xbit_r41_c142 bl_142 br_142 wl_41 vdd gnd cell_6t
Xbit_r42_c142 bl_142 br_142 wl_42 vdd gnd cell_6t
Xbit_r43_c142 bl_142 br_142 wl_43 vdd gnd cell_6t
Xbit_r44_c142 bl_142 br_142 wl_44 vdd gnd cell_6t
Xbit_r45_c142 bl_142 br_142 wl_45 vdd gnd cell_6t
Xbit_r46_c142 bl_142 br_142 wl_46 vdd gnd cell_6t
Xbit_r47_c142 bl_142 br_142 wl_47 vdd gnd cell_6t
Xbit_r48_c142 bl_142 br_142 wl_48 vdd gnd cell_6t
Xbit_r49_c142 bl_142 br_142 wl_49 vdd gnd cell_6t
Xbit_r50_c142 bl_142 br_142 wl_50 vdd gnd cell_6t
Xbit_r51_c142 bl_142 br_142 wl_51 vdd gnd cell_6t
Xbit_r52_c142 bl_142 br_142 wl_52 vdd gnd cell_6t
Xbit_r53_c142 bl_142 br_142 wl_53 vdd gnd cell_6t
Xbit_r54_c142 bl_142 br_142 wl_54 vdd gnd cell_6t
Xbit_r55_c142 bl_142 br_142 wl_55 vdd gnd cell_6t
Xbit_r56_c142 bl_142 br_142 wl_56 vdd gnd cell_6t
Xbit_r57_c142 bl_142 br_142 wl_57 vdd gnd cell_6t
Xbit_r58_c142 bl_142 br_142 wl_58 vdd gnd cell_6t
Xbit_r59_c142 bl_142 br_142 wl_59 vdd gnd cell_6t
Xbit_r60_c142 bl_142 br_142 wl_60 vdd gnd cell_6t
Xbit_r61_c142 bl_142 br_142 wl_61 vdd gnd cell_6t
Xbit_r62_c142 bl_142 br_142 wl_62 vdd gnd cell_6t
Xbit_r63_c142 bl_142 br_142 wl_63 vdd gnd cell_6t
Xbit_r64_c142 bl_142 br_142 wl_64 vdd gnd cell_6t
Xbit_r65_c142 bl_142 br_142 wl_65 vdd gnd cell_6t
Xbit_r66_c142 bl_142 br_142 wl_66 vdd gnd cell_6t
Xbit_r67_c142 bl_142 br_142 wl_67 vdd gnd cell_6t
Xbit_r68_c142 bl_142 br_142 wl_68 vdd gnd cell_6t
Xbit_r69_c142 bl_142 br_142 wl_69 vdd gnd cell_6t
Xbit_r70_c142 bl_142 br_142 wl_70 vdd gnd cell_6t
Xbit_r71_c142 bl_142 br_142 wl_71 vdd gnd cell_6t
Xbit_r72_c142 bl_142 br_142 wl_72 vdd gnd cell_6t
Xbit_r73_c142 bl_142 br_142 wl_73 vdd gnd cell_6t
Xbit_r74_c142 bl_142 br_142 wl_74 vdd gnd cell_6t
Xbit_r75_c142 bl_142 br_142 wl_75 vdd gnd cell_6t
Xbit_r76_c142 bl_142 br_142 wl_76 vdd gnd cell_6t
Xbit_r77_c142 bl_142 br_142 wl_77 vdd gnd cell_6t
Xbit_r78_c142 bl_142 br_142 wl_78 vdd gnd cell_6t
Xbit_r79_c142 bl_142 br_142 wl_79 vdd gnd cell_6t
Xbit_r80_c142 bl_142 br_142 wl_80 vdd gnd cell_6t
Xbit_r81_c142 bl_142 br_142 wl_81 vdd gnd cell_6t
Xbit_r82_c142 bl_142 br_142 wl_82 vdd gnd cell_6t
Xbit_r83_c142 bl_142 br_142 wl_83 vdd gnd cell_6t
Xbit_r84_c142 bl_142 br_142 wl_84 vdd gnd cell_6t
Xbit_r85_c142 bl_142 br_142 wl_85 vdd gnd cell_6t
Xbit_r86_c142 bl_142 br_142 wl_86 vdd gnd cell_6t
Xbit_r87_c142 bl_142 br_142 wl_87 vdd gnd cell_6t
Xbit_r88_c142 bl_142 br_142 wl_88 vdd gnd cell_6t
Xbit_r89_c142 bl_142 br_142 wl_89 vdd gnd cell_6t
Xbit_r90_c142 bl_142 br_142 wl_90 vdd gnd cell_6t
Xbit_r91_c142 bl_142 br_142 wl_91 vdd gnd cell_6t
Xbit_r92_c142 bl_142 br_142 wl_92 vdd gnd cell_6t
Xbit_r93_c142 bl_142 br_142 wl_93 vdd gnd cell_6t
Xbit_r94_c142 bl_142 br_142 wl_94 vdd gnd cell_6t
Xbit_r95_c142 bl_142 br_142 wl_95 vdd gnd cell_6t
Xbit_r96_c142 bl_142 br_142 wl_96 vdd gnd cell_6t
Xbit_r97_c142 bl_142 br_142 wl_97 vdd gnd cell_6t
Xbit_r98_c142 bl_142 br_142 wl_98 vdd gnd cell_6t
Xbit_r99_c142 bl_142 br_142 wl_99 vdd gnd cell_6t
Xbit_r100_c142 bl_142 br_142 wl_100 vdd gnd cell_6t
Xbit_r101_c142 bl_142 br_142 wl_101 vdd gnd cell_6t
Xbit_r102_c142 bl_142 br_142 wl_102 vdd gnd cell_6t
Xbit_r103_c142 bl_142 br_142 wl_103 vdd gnd cell_6t
Xbit_r104_c142 bl_142 br_142 wl_104 vdd gnd cell_6t
Xbit_r105_c142 bl_142 br_142 wl_105 vdd gnd cell_6t
Xbit_r106_c142 bl_142 br_142 wl_106 vdd gnd cell_6t
Xbit_r107_c142 bl_142 br_142 wl_107 vdd gnd cell_6t
Xbit_r108_c142 bl_142 br_142 wl_108 vdd gnd cell_6t
Xbit_r109_c142 bl_142 br_142 wl_109 vdd gnd cell_6t
Xbit_r110_c142 bl_142 br_142 wl_110 vdd gnd cell_6t
Xbit_r111_c142 bl_142 br_142 wl_111 vdd gnd cell_6t
Xbit_r112_c142 bl_142 br_142 wl_112 vdd gnd cell_6t
Xbit_r113_c142 bl_142 br_142 wl_113 vdd gnd cell_6t
Xbit_r114_c142 bl_142 br_142 wl_114 vdd gnd cell_6t
Xbit_r115_c142 bl_142 br_142 wl_115 vdd gnd cell_6t
Xbit_r116_c142 bl_142 br_142 wl_116 vdd gnd cell_6t
Xbit_r117_c142 bl_142 br_142 wl_117 vdd gnd cell_6t
Xbit_r118_c142 bl_142 br_142 wl_118 vdd gnd cell_6t
Xbit_r119_c142 bl_142 br_142 wl_119 vdd gnd cell_6t
Xbit_r120_c142 bl_142 br_142 wl_120 vdd gnd cell_6t
Xbit_r121_c142 bl_142 br_142 wl_121 vdd gnd cell_6t
Xbit_r122_c142 bl_142 br_142 wl_122 vdd gnd cell_6t
Xbit_r123_c142 bl_142 br_142 wl_123 vdd gnd cell_6t
Xbit_r124_c142 bl_142 br_142 wl_124 vdd gnd cell_6t
Xbit_r125_c142 bl_142 br_142 wl_125 vdd gnd cell_6t
Xbit_r126_c142 bl_142 br_142 wl_126 vdd gnd cell_6t
Xbit_r127_c142 bl_142 br_142 wl_127 vdd gnd cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd cell_6t
Xbit_r1_c143 bl_143 br_143 wl_1 vdd gnd cell_6t
Xbit_r2_c143 bl_143 br_143 wl_2 vdd gnd cell_6t
Xbit_r3_c143 bl_143 br_143 wl_3 vdd gnd cell_6t
Xbit_r4_c143 bl_143 br_143 wl_4 vdd gnd cell_6t
Xbit_r5_c143 bl_143 br_143 wl_5 vdd gnd cell_6t
Xbit_r6_c143 bl_143 br_143 wl_6 vdd gnd cell_6t
Xbit_r7_c143 bl_143 br_143 wl_7 vdd gnd cell_6t
Xbit_r8_c143 bl_143 br_143 wl_8 vdd gnd cell_6t
Xbit_r9_c143 bl_143 br_143 wl_9 vdd gnd cell_6t
Xbit_r10_c143 bl_143 br_143 wl_10 vdd gnd cell_6t
Xbit_r11_c143 bl_143 br_143 wl_11 vdd gnd cell_6t
Xbit_r12_c143 bl_143 br_143 wl_12 vdd gnd cell_6t
Xbit_r13_c143 bl_143 br_143 wl_13 vdd gnd cell_6t
Xbit_r14_c143 bl_143 br_143 wl_14 vdd gnd cell_6t
Xbit_r15_c143 bl_143 br_143 wl_15 vdd gnd cell_6t
Xbit_r16_c143 bl_143 br_143 wl_16 vdd gnd cell_6t
Xbit_r17_c143 bl_143 br_143 wl_17 vdd gnd cell_6t
Xbit_r18_c143 bl_143 br_143 wl_18 vdd gnd cell_6t
Xbit_r19_c143 bl_143 br_143 wl_19 vdd gnd cell_6t
Xbit_r20_c143 bl_143 br_143 wl_20 vdd gnd cell_6t
Xbit_r21_c143 bl_143 br_143 wl_21 vdd gnd cell_6t
Xbit_r22_c143 bl_143 br_143 wl_22 vdd gnd cell_6t
Xbit_r23_c143 bl_143 br_143 wl_23 vdd gnd cell_6t
Xbit_r24_c143 bl_143 br_143 wl_24 vdd gnd cell_6t
Xbit_r25_c143 bl_143 br_143 wl_25 vdd gnd cell_6t
Xbit_r26_c143 bl_143 br_143 wl_26 vdd gnd cell_6t
Xbit_r27_c143 bl_143 br_143 wl_27 vdd gnd cell_6t
Xbit_r28_c143 bl_143 br_143 wl_28 vdd gnd cell_6t
Xbit_r29_c143 bl_143 br_143 wl_29 vdd gnd cell_6t
Xbit_r30_c143 bl_143 br_143 wl_30 vdd gnd cell_6t
Xbit_r31_c143 bl_143 br_143 wl_31 vdd gnd cell_6t
Xbit_r32_c143 bl_143 br_143 wl_32 vdd gnd cell_6t
Xbit_r33_c143 bl_143 br_143 wl_33 vdd gnd cell_6t
Xbit_r34_c143 bl_143 br_143 wl_34 vdd gnd cell_6t
Xbit_r35_c143 bl_143 br_143 wl_35 vdd gnd cell_6t
Xbit_r36_c143 bl_143 br_143 wl_36 vdd gnd cell_6t
Xbit_r37_c143 bl_143 br_143 wl_37 vdd gnd cell_6t
Xbit_r38_c143 bl_143 br_143 wl_38 vdd gnd cell_6t
Xbit_r39_c143 bl_143 br_143 wl_39 vdd gnd cell_6t
Xbit_r40_c143 bl_143 br_143 wl_40 vdd gnd cell_6t
Xbit_r41_c143 bl_143 br_143 wl_41 vdd gnd cell_6t
Xbit_r42_c143 bl_143 br_143 wl_42 vdd gnd cell_6t
Xbit_r43_c143 bl_143 br_143 wl_43 vdd gnd cell_6t
Xbit_r44_c143 bl_143 br_143 wl_44 vdd gnd cell_6t
Xbit_r45_c143 bl_143 br_143 wl_45 vdd gnd cell_6t
Xbit_r46_c143 bl_143 br_143 wl_46 vdd gnd cell_6t
Xbit_r47_c143 bl_143 br_143 wl_47 vdd gnd cell_6t
Xbit_r48_c143 bl_143 br_143 wl_48 vdd gnd cell_6t
Xbit_r49_c143 bl_143 br_143 wl_49 vdd gnd cell_6t
Xbit_r50_c143 bl_143 br_143 wl_50 vdd gnd cell_6t
Xbit_r51_c143 bl_143 br_143 wl_51 vdd gnd cell_6t
Xbit_r52_c143 bl_143 br_143 wl_52 vdd gnd cell_6t
Xbit_r53_c143 bl_143 br_143 wl_53 vdd gnd cell_6t
Xbit_r54_c143 bl_143 br_143 wl_54 vdd gnd cell_6t
Xbit_r55_c143 bl_143 br_143 wl_55 vdd gnd cell_6t
Xbit_r56_c143 bl_143 br_143 wl_56 vdd gnd cell_6t
Xbit_r57_c143 bl_143 br_143 wl_57 vdd gnd cell_6t
Xbit_r58_c143 bl_143 br_143 wl_58 vdd gnd cell_6t
Xbit_r59_c143 bl_143 br_143 wl_59 vdd gnd cell_6t
Xbit_r60_c143 bl_143 br_143 wl_60 vdd gnd cell_6t
Xbit_r61_c143 bl_143 br_143 wl_61 vdd gnd cell_6t
Xbit_r62_c143 bl_143 br_143 wl_62 vdd gnd cell_6t
Xbit_r63_c143 bl_143 br_143 wl_63 vdd gnd cell_6t
Xbit_r64_c143 bl_143 br_143 wl_64 vdd gnd cell_6t
Xbit_r65_c143 bl_143 br_143 wl_65 vdd gnd cell_6t
Xbit_r66_c143 bl_143 br_143 wl_66 vdd gnd cell_6t
Xbit_r67_c143 bl_143 br_143 wl_67 vdd gnd cell_6t
Xbit_r68_c143 bl_143 br_143 wl_68 vdd gnd cell_6t
Xbit_r69_c143 bl_143 br_143 wl_69 vdd gnd cell_6t
Xbit_r70_c143 bl_143 br_143 wl_70 vdd gnd cell_6t
Xbit_r71_c143 bl_143 br_143 wl_71 vdd gnd cell_6t
Xbit_r72_c143 bl_143 br_143 wl_72 vdd gnd cell_6t
Xbit_r73_c143 bl_143 br_143 wl_73 vdd gnd cell_6t
Xbit_r74_c143 bl_143 br_143 wl_74 vdd gnd cell_6t
Xbit_r75_c143 bl_143 br_143 wl_75 vdd gnd cell_6t
Xbit_r76_c143 bl_143 br_143 wl_76 vdd gnd cell_6t
Xbit_r77_c143 bl_143 br_143 wl_77 vdd gnd cell_6t
Xbit_r78_c143 bl_143 br_143 wl_78 vdd gnd cell_6t
Xbit_r79_c143 bl_143 br_143 wl_79 vdd gnd cell_6t
Xbit_r80_c143 bl_143 br_143 wl_80 vdd gnd cell_6t
Xbit_r81_c143 bl_143 br_143 wl_81 vdd gnd cell_6t
Xbit_r82_c143 bl_143 br_143 wl_82 vdd gnd cell_6t
Xbit_r83_c143 bl_143 br_143 wl_83 vdd gnd cell_6t
Xbit_r84_c143 bl_143 br_143 wl_84 vdd gnd cell_6t
Xbit_r85_c143 bl_143 br_143 wl_85 vdd gnd cell_6t
Xbit_r86_c143 bl_143 br_143 wl_86 vdd gnd cell_6t
Xbit_r87_c143 bl_143 br_143 wl_87 vdd gnd cell_6t
Xbit_r88_c143 bl_143 br_143 wl_88 vdd gnd cell_6t
Xbit_r89_c143 bl_143 br_143 wl_89 vdd gnd cell_6t
Xbit_r90_c143 bl_143 br_143 wl_90 vdd gnd cell_6t
Xbit_r91_c143 bl_143 br_143 wl_91 vdd gnd cell_6t
Xbit_r92_c143 bl_143 br_143 wl_92 vdd gnd cell_6t
Xbit_r93_c143 bl_143 br_143 wl_93 vdd gnd cell_6t
Xbit_r94_c143 bl_143 br_143 wl_94 vdd gnd cell_6t
Xbit_r95_c143 bl_143 br_143 wl_95 vdd gnd cell_6t
Xbit_r96_c143 bl_143 br_143 wl_96 vdd gnd cell_6t
Xbit_r97_c143 bl_143 br_143 wl_97 vdd gnd cell_6t
Xbit_r98_c143 bl_143 br_143 wl_98 vdd gnd cell_6t
Xbit_r99_c143 bl_143 br_143 wl_99 vdd gnd cell_6t
Xbit_r100_c143 bl_143 br_143 wl_100 vdd gnd cell_6t
Xbit_r101_c143 bl_143 br_143 wl_101 vdd gnd cell_6t
Xbit_r102_c143 bl_143 br_143 wl_102 vdd gnd cell_6t
Xbit_r103_c143 bl_143 br_143 wl_103 vdd gnd cell_6t
Xbit_r104_c143 bl_143 br_143 wl_104 vdd gnd cell_6t
Xbit_r105_c143 bl_143 br_143 wl_105 vdd gnd cell_6t
Xbit_r106_c143 bl_143 br_143 wl_106 vdd gnd cell_6t
Xbit_r107_c143 bl_143 br_143 wl_107 vdd gnd cell_6t
Xbit_r108_c143 bl_143 br_143 wl_108 vdd gnd cell_6t
Xbit_r109_c143 bl_143 br_143 wl_109 vdd gnd cell_6t
Xbit_r110_c143 bl_143 br_143 wl_110 vdd gnd cell_6t
Xbit_r111_c143 bl_143 br_143 wl_111 vdd gnd cell_6t
Xbit_r112_c143 bl_143 br_143 wl_112 vdd gnd cell_6t
Xbit_r113_c143 bl_143 br_143 wl_113 vdd gnd cell_6t
Xbit_r114_c143 bl_143 br_143 wl_114 vdd gnd cell_6t
Xbit_r115_c143 bl_143 br_143 wl_115 vdd gnd cell_6t
Xbit_r116_c143 bl_143 br_143 wl_116 vdd gnd cell_6t
Xbit_r117_c143 bl_143 br_143 wl_117 vdd gnd cell_6t
Xbit_r118_c143 bl_143 br_143 wl_118 vdd gnd cell_6t
Xbit_r119_c143 bl_143 br_143 wl_119 vdd gnd cell_6t
Xbit_r120_c143 bl_143 br_143 wl_120 vdd gnd cell_6t
Xbit_r121_c143 bl_143 br_143 wl_121 vdd gnd cell_6t
Xbit_r122_c143 bl_143 br_143 wl_122 vdd gnd cell_6t
Xbit_r123_c143 bl_143 br_143 wl_123 vdd gnd cell_6t
Xbit_r124_c143 bl_143 br_143 wl_124 vdd gnd cell_6t
Xbit_r125_c143 bl_143 br_143 wl_125 vdd gnd cell_6t
Xbit_r126_c143 bl_143 br_143 wl_126 vdd gnd cell_6t
Xbit_r127_c143 bl_143 br_143 wl_127 vdd gnd cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd cell_6t
Xbit_r1_c144 bl_144 br_144 wl_1 vdd gnd cell_6t
Xbit_r2_c144 bl_144 br_144 wl_2 vdd gnd cell_6t
Xbit_r3_c144 bl_144 br_144 wl_3 vdd gnd cell_6t
Xbit_r4_c144 bl_144 br_144 wl_4 vdd gnd cell_6t
Xbit_r5_c144 bl_144 br_144 wl_5 vdd gnd cell_6t
Xbit_r6_c144 bl_144 br_144 wl_6 vdd gnd cell_6t
Xbit_r7_c144 bl_144 br_144 wl_7 vdd gnd cell_6t
Xbit_r8_c144 bl_144 br_144 wl_8 vdd gnd cell_6t
Xbit_r9_c144 bl_144 br_144 wl_9 vdd gnd cell_6t
Xbit_r10_c144 bl_144 br_144 wl_10 vdd gnd cell_6t
Xbit_r11_c144 bl_144 br_144 wl_11 vdd gnd cell_6t
Xbit_r12_c144 bl_144 br_144 wl_12 vdd gnd cell_6t
Xbit_r13_c144 bl_144 br_144 wl_13 vdd gnd cell_6t
Xbit_r14_c144 bl_144 br_144 wl_14 vdd gnd cell_6t
Xbit_r15_c144 bl_144 br_144 wl_15 vdd gnd cell_6t
Xbit_r16_c144 bl_144 br_144 wl_16 vdd gnd cell_6t
Xbit_r17_c144 bl_144 br_144 wl_17 vdd gnd cell_6t
Xbit_r18_c144 bl_144 br_144 wl_18 vdd gnd cell_6t
Xbit_r19_c144 bl_144 br_144 wl_19 vdd gnd cell_6t
Xbit_r20_c144 bl_144 br_144 wl_20 vdd gnd cell_6t
Xbit_r21_c144 bl_144 br_144 wl_21 vdd gnd cell_6t
Xbit_r22_c144 bl_144 br_144 wl_22 vdd gnd cell_6t
Xbit_r23_c144 bl_144 br_144 wl_23 vdd gnd cell_6t
Xbit_r24_c144 bl_144 br_144 wl_24 vdd gnd cell_6t
Xbit_r25_c144 bl_144 br_144 wl_25 vdd gnd cell_6t
Xbit_r26_c144 bl_144 br_144 wl_26 vdd gnd cell_6t
Xbit_r27_c144 bl_144 br_144 wl_27 vdd gnd cell_6t
Xbit_r28_c144 bl_144 br_144 wl_28 vdd gnd cell_6t
Xbit_r29_c144 bl_144 br_144 wl_29 vdd gnd cell_6t
Xbit_r30_c144 bl_144 br_144 wl_30 vdd gnd cell_6t
Xbit_r31_c144 bl_144 br_144 wl_31 vdd gnd cell_6t
Xbit_r32_c144 bl_144 br_144 wl_32 vdd gnd cell_6t
Xbit_r33_c144 bl_144 br_144 wl_33 vdd gnd cell_6t
Xbit_r34_c144 bl_144 br_144 wl_34 vdd gnd cell_6t
Xbit_r35_c144 bl_144 br_144 wl_35 vdd gnd cell_6t
Xbit_r36_c144 bl_144 br_144 wl_36 vdd gnd cell_6t
Xbit_r37_c144 bl_144 br_144 wl_37 vdd gnd cell_6t
Xbit_r38_c144 bl_144 br_144 wl_38 vdd gnd cell_6t
Xbit_r39_c144 bl_144 br_144 wl_39 vdd gnd cell_6t
Xbit_r40_c144 bl_144 br_144 wl_40 vdd gnd cell_6t
Xbit_r41_c144 bl_144 br_144 wl_41 vdd gnd cell_6t
Xbit_r42_c144 bl_144 br_144 wl_42 vdd gnd cell_6t
Xbit_r43_c144 bl_144 br_144 wl_43 vdd gnd cell_6t
Xbit_r44_c144 bl_144 br_144 wl_44 vdd gnd cell_6t
Xbit_r45_c144 bl_144 br_144 wl_45 vdd gnd cell_6t
Xbit_r46_c144 bl_144 br_144 wl_46 vdd gnd cell_6t
Xbit_r47_c144 bl_144 br_144 wl_47 vdd gnd cell_6t
Xbit_r48_c144 bl_144 br_144 wl_48 vdd gnd cell_6t
Xbit_r49_c144 bl_144 br_144 wl_49 vdd gnd cell_6t
Xbit_r50_c144 bl_144 br_144 wl_50 vdd gnd cell_6t
Xbit_r51_c144 bl_144 br_144 wl_51 vdd gnd cell_6t
Xbit_r52_c144 bl_144 br_144 wl_52 vdd gnd cell_6t
Xbit_r53_c144 bl_144 br_144 wl_53 vdd gnd cell_6t
Xbit_r54_c144 bl_144 br_144 wl_54 vdd gnd cell_6t
Xbit_r55_c144 bl_144 br_144 wl_55 vdd gnd cell_6t
Xbit_r56_c144 bl_144 br_144 wl_56 vdd gnd cell_6t
Xbit_r57_c144 bl_144 br_144 wl_57 vdd gnd cell_6t
Xbit_r58_c144 bl_144 br_144 wl_58 vdd gnd cell_6t
Xbit_r59_c144 bl_144 br_144 wl_59 vdd gnd cell_6t
Xbit_r60_c144 bl_144 br_144 wl_60 vdd gnd cell_6t
Xbit_r61_c144 bl_144 br_144 wl_61 vdd gnd cell_6t
Xbit_r62_c144 bl_144 br_144 wl_62 vdd gnd cell_6t
Xbit_r63_c144 bl_144 br_144 wl_63 vdd gnd cell_6t
Xbit_r64_c144 bl_144 br_144 wl_64 vdd gnd cell_6t
Xbit_r65_c144 bl_144 br_144 wl_65 vdd gnd cell_6t
Xbit_r66_c144 bl_144 br_144 wl_66 vdd gnd cell_6t
Xbit_r67_c144 bl_144 br_144 wl_67 vdd gnd cell_6t
Xbit_r68_c144 bl_144 br_144 wl_68 vdd gnd cell_6t
Xbit_r69_c144 bl_144 br_144 wl_69 vdd gnd cell_6t
Xbit_r70_c144 bl_144 br_144 wl_70 vdd gnd cell_6t
Xbit_r71_c144 bl_144 br_144 wl_71 vdd gnd cell_6t
Xbit_r72_c144 bl_144 br_144 wl_72 vdd gnd cell_6t
Xbit_r73_c144 bl_144 br_144 wl_73 vdd gnd cell_6t
Xbit_r74_c144 bl_144 br_144 wl_74 vdd gnd cell_6t
Xbit_r75_c144 bl_144 br_144 wl_75 vdd gnd cell_6t
Xbit_r76_c144 bl_144 br_144 wl_76 vdd gnd cell_6t
Xbit_r77_c144 bl_144 br_144 wl_77 vdd gnd cell_6t
Xbit_r78_c144 bl_144 br_144 wl_78 vdd gnd cell_6t
Xbit_r79_c144 bl_144 br_144 wl_79 vdd gnd cell_6t
Xbit_r80_c144 bl_144 br_144 wl_80 vdd gnd cell_6t
Xbit_r81_c144 bl_144 br_144 wl_81 vdd gnd cell_6t
Xbit_r82_c144 bl_144 br_144 wl_82 vdd gnd cell_6t
Xbit_r83_c144 bl_144 br_144 wl_83 vdd gnd cell_6t
Xbit_r84_c144 bl_144 br_144 wl_84 vdd gnd cell_6t
Xbit_r85_c144 bl_144 br_144 wl_85 vdd gnd cell_6t
Xbit_r86_c144 bl_144 br_144 wl_86 vdd gnd cell_6t
Xbit_r87_c144 bl_144 br_144 wl_87 vdd gnd cell_6t
Xbit_r88_c144 bl_144 br_144 wl_88 vdd gnd cell_6t
Xbit_r89_c144 bl_144 br_144 wl_89 vdd gnd cell_6t
Xbit_r90_c144 bl_144 br_144 wl_90 vdd gnd cell_6t
Xbit_r91_c144 bl_144 br_144 wl_91 vdd gnd cell_6t
Xbit_r92_c144 bl_144 br_144 wl_92 vdd gnd cell_6t
Xbit_r93_c144 bl_144 br_144 wl_93 vdd gnd cell_6t
Xbit_r94_c144 bl_144 br_144 wl_94 vdd gnd cell_6t
Xbit_r95_c144 bl_144 br_144 wl_95 vdd gnd cell_6t
Xbit_r96_c144 bl_144 br_144 wl_96 vdd gnd cell_6t
Xbit_r97_c144 bl_144 br_144 wl_97 vdd gnd cell_6t
Xbit_r98_c144 bl_144 br_144 wl_98 vdd gnd cell_6t
Xbit_r99_c144 bl_144 br_144 wl_99 vdd gnd cell_6t
Xbit_r100_c144 bl_144 br_144 wl_100 vdd gnd cell_6t
Xbit_r101_c144 bl_144 br_144 wl_101 vdd gnd cell_6t
Xbit_r102_c144 bl_144 br_144 wl_102 vdd gnd cell_6t
Xbit_r103_c144 bl_144 br_144 wl_103 vdd gnd cell_6t
Xbit_r104_c144 bl_144 br_144 wl_104 vdd gnd cell_6t
Xbit_r105_c144 bl_144 br_144 wl_105 vdd gnd cell_6t
Xbit_r106_c144 bl_144 br_144 wl_106 vdd gnd cell_6t
Xbit_r107_c144 bl_144 br_144 wl_107 vdd gnd cell_6t
Xbit_r108_c144 bl_144 br_144 wl_108 vdd gnd cell_6t
Xbit_r109_c144 bl_144 br_144 wl_109 vdd gnd cell_6t
Xbit_r110_c144 bl_144 br_144 wl_110 vdd gnd cell_6t
Xbit_r111_c144 bl_144 br_144 wl_111 vdd gnd cell_6t
Xbit_r112_c144 bl_144 br_144 wl_112 vdd gnd cell_6t
Xbit_r113_c144 bl_144 br_144 wl_113 vdd gnd cell_6t
Xbit_r114_c144 bl_144 br_144 wl_114 vdd gnd cell_6t
Xbit_r115_c144 bl_144 br_144 wl_115 vdd gnd cell_6t
Xbit_r116_c144 bl_144 br_144 wl_116 vdd gnd cell_6t
Xbit_r117_c144 bl_144 br_144 wl_117 vdd gnd cell_6t
Xbit_r118_c144 bl_144 br_144 wl_118 vdd gnd cell_6t
Xbit_r119_c144 bl_144 br_144 wl_119 vdd gnd cell_6t
Xbit_r120_c144 bl_144 br_144 wl_120 vdd gnd cell_6t
Xbit_r121_c144 bl_144 br_144 wl_121 vdd gnd cell_6t
Xbit_r122_c144 bl_144 br_144 wl_122 vdd gnd cell_6t
Xbit_r123_c144 bl_144 br_144 wl_123 vdd gnd cell_6t
Xbit_r124_c144 bl_144 br_144 wl_124 vdd gnd cell_6t
Xbit_r125_c144 bl_144 br_144 wl_125 vdd gnd cell_6t
Xbit_r126_c144 bl_144 br_144 wl_126 vdd gnd cell_6t
Xbit_r127_c144 bl_144 br_144 wl_127 vdd gnd cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd cell_6t
Xbit_r1_c145 bl_145 br_145 wl_1 vdd gnd cell_6t
Xbit_r2_c145 bl_145 br_145 wl_2 vdd gnd cell_6t
Xbit_r3_c145 bl_145 br_145 wl_3 vdd gnd cell_6t
Xbit_r4_c145 bl_145 br_145 wl_4 vdd gnd cell_6t
Xbit_r5_c145 bl_145 br_145 wl_5 vdd gnd cell_6t
Xbit_r6_c145 bl_145 br_145 wl_6 vdd gnd cell_6t
Xbit_r7_c145 bl_145 br_145 wl_7 vdd gnd cell_6t
Xbit_r8_c145 bl_145 br_145 wl_8 vdd gnd cell_6t
Xbit_r9_c145 bl_145 br_145 wl_9 vdd gnd cell_6t
Xbit_r10_c145 bl_145 br_145 wl_10 vdd gnd cell_6t
Xbit_r11_c145 bl_145 br_145 wl_11 vdd gnd cell_6t
Xbit_r12_c145 bl_145 br_145 wl_12 vdd gnd cell_6t
Xbit_r13_c145 bl_145 br_145 wl_13 vdd gnd cell_6t
Xbit_r14_c145 bl_145 br_145 wl_14 vdd gnd cell_6t
Xbit_r15_c145 bl_145 br_145 wl_15 vdd gnd cell_6t
Xbit_r16_c145 bl_145 br_145 wl_16 vdd gnd cell_6t
Xbit_r17_c145 bl_145 br_145 wl_17 vdd gnd cell_6t
Xbit_r18_c145 bl_145 br_145 wl_18 vdd gnd cell_6t
Xbit_r19_c145 bl_145 br_145 wl_19 vdd gnd cell_6t
Xbit_r20_c145 bl_145 br_145 wl_20 vdd gnd cell_6t
Xbit_r21_c145 bl_145 br_145 wl_21 vdd gnd cell_6t
Xbit_r22_c145 bl_145 br_145 wl_22 vdd gnd cell_6t
Xbit_r23_c145 bl_145 br_145 wl_23 vdd gnd cell_6t
Xbit_r24_c145 bl_145 br_145 wl_24 vdd gnd cell_6t
Xbit_r25_c145 bl_145 br_145 wl_25 vdd gnd cell_6t
Xbit_r26_c145 bl_145 br_145 wl_26 vdd gnd cell_6t
Xbit_r27_c145 bl_145 br_145 wl_27 vdd gnd cell_6t
Xbit_r28_c145 bl_145 br_145 wl_28 vdd gnd cell_6t
Xbit_r29_c145 bl_145 br_145 wl_29 vdd gnd cell_6t
Xbit_r30_c145 bl_145 br_145 wl_30 vdd gnd cell_6t
Xbit_r31_c145 bl_145 br_145 wl_31 vdd gnd cell_6t
Xbit_r32_c145 bl_145 br_145 wl_32 vdd gnd cell_6t
Xbit_r33_c145 bl_145 br_145 wl_33 vdd gnd cell_6t
Xbit_r34_c145 bl_145 br_145 wl_34 vdd gnd cell_6t
Xbit_r35_c145 bl_145 br_145 wl_35 vdd gnd cell_6t
Xbit_r36_c145 bl_145 br_145 wl_36 vdd gnd cell_6t
Xbit_r37_c145 bl_145 br_145 wl_37 vdd gnd cell_6t
Xbit_r38_c145 bl_145 br_145 wl_38 vdd gnd cell_6t
Xbit_r39_c145 bl_145 br_145 wl_39 vdd gnd cell_6t
Xbit_r40_c145 bl_145 br_145 wl_40 vdd gnd cell_6t
Xbit_r41_c145 bl_145 br_145 wl_41 vdd gnd cell_6t
Xbit_r42_c145 bl_145 br_145 wl_42 vdd gnd cell_6t
Xbit_r43_c145 bl_145 br_145 wl_43 vdd gnd cell_6t
Xbit_r44_c145 bl_145 br_145 wl_44 vdd gnd cell_6t
Xbit_r45_c145 bl_145 br_145 wl_45 vdd gnd cell_6t
Xbit_r46_c145 bl_145 br_145 wl_46 vdd gnd cell_6t
Xbit_r47_c145 bl_145 br_145 wl_47 vdd gnd cell_6t
Xbit_r48_c145 bl_145 br_145 wl_48 vdd gnd cell_6t
Xbit_r49_c145 bl_145 br_145 wl_49 vdd gnd cell_6t
Xbit_r50_c145 bl_145 br_145 wl_50 vdd gnd cell_6t
Xbit_r51_c145 bl_145 br_145 wl_51 vdd gnd cell_6t
Xbit_r52_c145 bl_145 br_145 wl_52 vdd gnd cell_6t
Xbit_r53_c145 bl_145 br_145 wl_53 vdd gnd cell_6t
Xbit_r54_c145 bl_145 br_145 wl_54 vdd gnd cell_6t
Xbit_r55_c145 bl_145 br_145 wl_55 vdd gnd cell_6t
Xbit_r56_c145 bl_145 br_145 wl_56 vdd gnd cell_6t
Xbit_r57_c145 bl_145 br_145 wl_57 vdd gnd cell_6t
Xbit_r58_c145 bl_145 br_145 wl_58 vdd gnd cell_6t
Xbit_r59_c145 bl_145 br_145 wl_59 vdd gnd cell_6t
Xbit_r60_c145 bl_145 br_145 wl_60 vdd gnd cell_6t
Xbit_r61_c145 bl_145 br_145 wl_61 vdd gnd cell_6t
Xbit_r62_c145 bl_145 br_145 wl_62 vdd gnd cell_6t
Xbit_r63_c145 bl_145 br_145 wl_63 vdd gnd cell_6t
Xbit_r64_c145 bl_145 br_145 wl_64 vdd gnd cell_6t
Xbit_r65_c145 bl_145 br_145 wl_65 vdd gnd cell_6t
Xbit_r66_c145 bl_145 br_145 wl_66 vdd gnd cell_6t
Xbit_r67_c145 bl_145 br_145 wl_67 vdd gnd cell_6t
Xbit_r68_c145 bl_145 br_145 wl_68 vdd gnd cell_6t
Xbit_r69_c145 bl_145 br_145 wl_69 vdd gnd cell_6t
Xbit_r70_c145 bl_145 br_145 wl_70 vdd gnd cell_6t
Xbit_r71_c145 bl_145 br_145 wl_71 vdd gnd cell_6t
Xbit_r72_c145 bl_145 br_145 wl_72 vdd gnd cell_6t
Xbit_r73_c145 bl_145 br_145 wl_73 vdd gnd cell_6t
Xbit_r74_c145 bl_145 br_145 wl_74 vdd gnd cell_6t
Xbit_r75_c145 bl_145 br_145 wl_75 vdd gnd cell_6t
Xbit_r76_c145 bl_145 br_145 wl_76 vdd gnd cell_6t
Xbit_r77_c145 bl_145 br_145 wl_77 vdd gnd cell_6t
Xbit_r78_c145 bl_145 br_145 wl_78 vdd gnd cell_6t
Xbit_r79_c145 bl_145 br_145 wl_79 vdd gnd cell_6t
Xbit_r80_c145 bl_145 br_145 wl_80 vdd gnd cell_6t
Xbit_r81_c145 bl_145 br_145 wl_81 vdd gnd cell_6t
Xbit_r82_c145 bl_145 br_145 wl_82 vdd gnd cell_6t
Xbit_r83_c145 bl_145 br_145 wl_83 vdd gnd cell_6t
Xbit_r84_c145 bl_145 br_145 wl_84 vdd gnd cell_6t
Xbit_r85_c145 bl_145 br_145 wl_85 vdd gnd cell_6t
Xbit_r86_c145 bl_145 br_145 wl_86 vdd gnd cell_6t
Xbit_r87_c145 bl_145 br_145 wl_87 vdd gnd cell_6t
Xbit_r88_c145 bl_145 br_145 wl_88 vdd gnd cell_6t
Xbit_r89_c145 bl_145 br_145 wl_89 vdd gnd cell_6t
Xbit_r90_c145 bl_145 br_145 wl_90 vdd gnd cell_6t
Xbit_r91_c145 bl_145 br_145 wl_91 vdd gnd cell_6t
Xbit_r92_c145 bl_145 br_145 wl_92 vdd gnd cell_6t
Xbit_r93_c145 bl_145 br_145 wl_93 vdd gnd cell_6t
Xbit_r94_c145 bl_145 br_145 wl_94 vdd gnd cell_6t
Xbit_r95_c145 bl_145 br_145 wl_95 vdd gnd cell_6t
Xbit_r96_c145 bl_145 br_145 wl_96 vdd gnd cell_6t
Xbit_r97_c145 bl_145 br_145 wl_97 vdd gnd cell_6t
Xbit_r98_c145 bl_145 br_145 wl_98 vdd gnd cell_6t
Xbit_r99_c145 bl_145 br_145 wl_99 vdd gnd cell_6t
Xbit_r100_c145 bl_145 br_145 wl_100 vdd gnd cell_6t
Xbit_r101_c145 bl_145 br_145 wl_101 vdd gnd cell_6t
Xbit_r102_c145 bl_145 br_145 wl_102 vdd gnd cell_6t
Xbit_r103_c145 bl_145 br_145 wl_103 vdd gnd cell_6t
Xbit_r104_c145 bl_145 br_145 wl_104 vdd gnd cell_6t
Xbit_r105_c145 bl_145 br_145 wl_105 vdd gnd cell_6t
Xbit_r106_c145 bl_145 br_145 wl_106 vdd gnd cell_6t
Xbit_r107_c145 bl_145 br_145 wl_107 vdd gnd cell_6t
Xbit_r108_c145 bl_145 br_145 wl_108 vdd gnd cell_6t
Xbit_r109_c145 bl_145 br_145 wl_109 vdd gnd cell_6t
Xbit_r110_c145 bl_145 br_145 wl_110 vdd gnd cell_6t
Xbit_r111_c145 bl_145 br_145 wl_111 vdd gnd cell_6t
Xbit_r112_c145 bl_145 br_145 wl_112 vdd gnd cell_6t
Xbit_r113_c145 bl_145 br_145 wl_113 vdd gnd cell_6t
Xbit_r114_c145 bl_145 br_145 wl_114 vdd gnd cell_6t
Xbit_r115_c145 bl_145 br_145 wl_115 vdd gnd cell_6t
Xbit_r116_c145 bl_145 br_145 wl_116 vdd gnd cell_6t
Xbit_r117_c145 bl_145 br_145 wl_117 vdd gnd cell_6t
Xbit_r118_c145 bl_145 br_145 wl_118 vdd gnd cell_6t
Xbit_r119_c145 bl_145 br_145 wl_119 vdd gnd cell_6t
Xbit_r120_c145 bl_145 br_145 wl_120 vdd gnd cell_6t
Xbit_r121_c145 bl_145 br_145 wl_121 vdd gnd cell_6t
Xbit_r122_c145 bl_145 br_145 wl_122 vdd gnd cell_6t
Xbit_r123_c145 bl_145 br_145 wl_123 vdd gnd cell_6t
Xbit_r124_c145 bl_145 br_145 wl_124 vdd gnd cell_6t
Xbit_r125_c145 bl_145 br_145 wl_125 vdd gnd cell_6t
Xbit_r126_c145 bl_145 br_145 wl_126 vdd gnd cell_6t
Xbit_r127_c145 bl_145 br_145 wl_127 vdd gnd cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd cell_6t
Xbit_r1_c146 bl_146 br_146 wl_1 vdd gnd cell_6t
Xbit_r2_c146 bl_146 br_146 wl_2 vdd gnd cell_6t
Xbit_r3_c146 bl_146 br_146 wl_3 vdd gnd cell_6t
Xbit_r4_c146 bl_146 br_146 wl_4 vdd gnd cell_6t
Xbit_r5_c146 bl_146 br_146 wl_5 vdd gnd cell_6t
Xbit_r6_c146 bl_146 br_146 wl_6 vdd gnd cell_6t
Xbit_r7_c146 bl_146 br_146 wl_7 vdd gnd cell_6t
Xbit_r8_c146 bl_146 br_146 wl_8 vdd gnd cell_6t
Xbit_r9_c146 bl_146 br_146 wl_9 vdd gnd cell_6t
Xbit_r10_c146 bl_146 br_146 wl_10 vdd gnd cell_6t
Xbit_r11_c146 bl_146 br_146 wl_11 vdd gnd cell_6t
Xbit_r12_c146 bl_146 br_146 wl_12 vdd gnd cell_6t
Xbit_r13_c146 bl_146 br_146 wl_13 vdd gnd cell_6t
Xbit_r14_c146 bl_146 br_146 wl_14 vdd gnd cell_6t
Xbit_r15_c146 bl_146 br_146 wl_15 vdd gnd cell_6t
Xbit_r16_c146 bl_146 br_146 wl_16 vdd gnd cell_6t
Xbit_r17_c146 bl_146 br_146 wl_17 vdd gnd cell_6t
Xbit_r18_c146 bl_146 br_146 wl_18 vdd gnd cell_6t
Xbit_r19_c146 bl_146 br_146 wl_19 vdd gnd cell_6t
Xbit_r20_c146 bl_146 br_146 wl_20 vdd gnd cell_6t
Xbit_r21_c146 bl_146 br_146 wl_21 vdd gnd cell_6t
Xbit_r22_c146 bl_146 br_146 wl_22 vdd gnd cell_6t
Xbit_r23_c146 bl_146 br_146 wl_23 vdd gnd cell_6t
Xbit_r24_c146 bl_146 br_146 wl_24 vdd gnd cell_6t
Xbit_r25_c146 bl_146 br_146 wl_25 vdd gnd cell_6t
Xbit_r26_c146 bl_146 br_146 wl_26 vdd gnd cell_6t
Xbit_r27_c146 bl_146 br_146 wl_27 vdd gnd cell_6t
Xbit_r28_c146 bl_146 br_146 wl_28 vdd gnd cell_6t
Xbit_r29_c146 bl_146 br_146 wl_29 vdd gnd cell_6t
Xbit_r30_c146 bl_146 br_146 wl_30 vdd gnd cell_6t
Xbit_r31_c146 bl_146 br_146 wl_31 vdd gnd cell_6t
Xbit_r32_c146 bl_146 br_146 wl_32 vdd gnd cell_6t
Xbit_r33_c146 bl_146 br_146 wl_33 vdd gnd cell_6t
Xbit_r34_c146 bl_146 br_146 wl_34 vdd gnd cell_6t
Xbit_r35_c146 bl_146 br_146 wl_35 vdd gnd cell_6t
Xbit_r36_c146 bl_146 br_146 wl_36 vdd gnd cell_6t
Xbit_r37_c146 bl_146 br_146 wl_37 vdd gnd cell_6t
Xbit_r38_c146 bl_146 br_146 wl_38 vdd gnd cell_6t
Xbit_r39_c146 bl_146 br_146 wl_39 vdd gnd cell_6t
Xbit_r40_c146 bl_146 br_146 wl_40 vdd gnd cell_6t
Xbit_r41_c146 bl_146 br_146 wl_41 vdd gnd cell_6t
Xbit_r42_c146 bl_146 br_146 wl_42 vdd gnd cell_6t
Xbit_r43_c146 bl_146 br_146 wl_43 vdd gnd cell_6t
Xbit_r44_c146 bl_146 br_146 wl_44 vdd gnd cell_6t
Xbit_r45_c146 bl_146 br_146 wl_45 vdd gnd cell_6t
Xbit_r46_c146 bl_146 br_146 wl_46 vdd gnd cell_6t
Xbit_r47_c146 bl_146 br_146 wl_47 vdd gnd cell_6t
Xbit_r48_c146 bl_146 br_146 wl_48 vdd gnd cell_6t
Xbit_r49_c146 bl_146 br_146 wl_49 vdd gnd cell_6t
Xbit_r50_c146 bl_146 br_146 wl_50 vdd gnd cell_6t
Xbit_r51_c146 bl_146 br_146 wl_51 vdd gnd cell_6t
Xbit_r52_c146 bl_146 br_146 wl_52 vdd gnd cell_6t
Xbit_r53_c146 bl_146 br_146 wl_53 vdd gnd cell_6t
Xbit_r54_c146 bl_146 br_146 wl_54 vdd gnd cell_6t
Xbit_r55_c146 bl_146 br_146 wl_55 vdd gnd cell_6t
Xbit_r56_c146 bl_146 br_146 wl_56 vdd gnd cell_6t
Xbit_r57_c146 bl_146 br_146 wl_57 vdd gnd cell_6t
Xbit_r58_c146 bl_146 br_146 wl_58 vdd gnd cell_6t
Xbit_r59_c146 bl_146 br_146 wl_59 vdd gnd cell_6t
Xbit_r60_c146 bl_146 br_146 wl_60 vdd gnd cell_6t
Xbit_r61_c146 bl_146 br_146 wl_61 vdd gnd cell_6t
Xbit_r62_c146 bl_146 br_146 wl_62 vdd gnd cell_6t
Xbit_r63_c146 bl_146 br_146 wl_63 vdd gnd cell_6t
Xbit_r64_c146 bl_146 br_146 wl_64 vdd gnd cell_6t
Xbit_r65_c146 bl_146 br_146 wl_65 vdd gnd cell_6t
Xbit_r66_c146 bl_146 br_146 wl_66 vdd gnd cell_6t
Xbit_r67_c146 bl_146 br_146 wl_67 vdd gnd cell_6t
Xbit_r68_c146 bl_146 br_146 wl_68 vdd gnd cell_6t
Xbit_r69_c146 bl_146 br_146 wl_69 vdd gnd cell_6t
Xbit_r70_c146 bl_146 br_146 wl_70 vdd gnd cell_6t
Xbit_r71_c146 bl_146 br_146 wl_71 vdd gnd cell_6t
Xbit_r72_c146 bl_146 br_146 wl_72 vdd gnd cell_6t
Xbit_r73_c146 bl_146 br_146 wl_73 vdd gnd cell_6t
Xbit_r74_c146 bl_146 br_146 wl_74 vdd gnd cell_6t
Xbit_r75_c146 bl_146 br_146 wl_75 vdd gnd cell_6t
Xbit_r76_c146 bl_146 br_146 wl_76 vdd gnd cell_6t
Xbit_r77_c146 bl_146 br_146 wl_77 vdd gnd cell_6t
Xbit_r78_c146 bl_146 br_146 wl_78 vdd gnd cell_6t
Xbit_r79_c146 bl_146 br_146 wl_79 vdd gnd cell_6t
Xbit_r80_c146 bl_146 br_146 wl_80 vdd gnd cell_6t
Xbit_r81_c146 bl_146 br_146 wl_81 vdd gnd cell_6t
Xbit_r82_c146 bl_146 br_146 wl_82 vdd gnd cell_6t
Xbit_r83_c146 bl_146 br_146 wl_83 vdd gnd cell_6t
Xbit_r84_c146 bl_146 br_146 wl_84 vdd gnd cell_6t
Xbit_r85_c146 bl_146 br_146 wl_85 vdd gnd cell_6t
Xbit_r86_c146 bl_146 br_146 wl_86 vdd gnd cell_6t
Xbit_r87_c146 bl_146 br_146 wl_87 vdd gnd cell_6t
Xbit_r88_c146 bl_146 br_146 wl_88 vdd gnd cell_6t
Xbit_r89_c146 bl_146 br_146 wl_89 vdd gnd cell_6t
Xbit_r90_c146 bl_146 br_146 wl_90 vdd gnd cell_6t
Xbit_r91_c146 bl_146 br_146 wl_91 vdd gnd cell_6t
Xbit_r92_c146 bl_146 br_146 wl_92 vdd gnd cell_6t
Xbit_r93_c146 bl_146 br_146 wl_93 vdd gnd cell_6t
Xbit_r94_c146 bl_146 br_146 wl_94 vdd gnd cell_6t
Xbit_r95_c146 bl_146 br_146 wl_95 vdd gnd cell_6t
Xbit_r96_c146 bl_146 br_146 wl_96 vdd gnd cell_6t
Xbit_r97_c146 bl_146 br_146 wl_97 vdd gnd cell_6t
Xbit_r98_c146 bl_146 br_146 wl_98 vdd gnd cell_6t
Xbit_r99_c146 bl_146 br_146 wl_99 vdd gnd cell_6t
Xbit_r100_c146 bl_146 br_146 wl_100 vdd gnd cell_6t
Xbit_r101_c146 bl_146 br_146 wl_101 vdd gnd cell_6t
Xbit_r102_c146 bl_146 br_146 wl_102 vdd gnd cell_6t
Xbit_r103_c146 bl_146 br_146 wl_103 vdd gnd cell_6t
Xbit_r104_c146 bl_146 br_146 wl_104 vdd gnd cell_6t
Xbit_r105_c146 bl_146 br_146 wl_105 vdd gnd cell_6t
Xbit_r106_c146 bl_146 br_146 wl_106 vdd gnd cell_6t
Xbit_r107_c146 bl_146 br_146 wl_107 vdd gnd cell_6t
Xbit_r108_c146 bl_146 br_146 wl_108 vdd gnd cell_6t
Xbit_r109_c146 bl_146 br_146 wl_109 vdd gnd cell_6t
Xbit_r110_c146 bl_146 br_146 wl_110 vdd gnd cell_6t
Xbit_r111_c146 bl_146 br_146 wl_111 vdd gnd cell_6t
Xbit_r112_c146 bl_146 br_146 wl_112 vdd gnd cell_6t
Xbit_r113_c146 bl_146 br_146 wl_113 vdd gnd cell_6t
Xbit_r114_c146 bl_146 br_146 wl_114 vdd gnd cell_6t
Xbit_r115_c146 bl_146 br_146 wl_115 vdd gnd cell_6t
Xbit_r116_c146 bl_146 br_146 wl_116 vdd gnd cell_6t
Xbit_r117_c146 bl_146 br_146 wl_117 vdd gnd cell_6t
Xbit_r118_c146 bl_146 br_146 wl_118 vdd gnd cell_6t
Xbit_r119_c146 bl_146 br_146 wl_119 vdd gnd cell_6t
Xbit_r120_c146 bl_146 br_146 wl_120 vdd gnd cell_6t
Xbit_r121_c146 bl_146 br_146 wl_121 vdd gnd cell_6t
Xbit_r122_c146 bl_146 br_146 wl_122 vdd gnd cell_6t
Xbit_r123_c146 bl_146 br_146 wl_123 vdd gnd cell_6t
Xbit_r124_c146 bl_146 br_146 wl_124 vdd gnd cell_6t
Xbit_r125_c146 bl_146 br_146 wl_125 vdd gnd cell_6t
Xbit_r126_c146 bl_146 br_146 wl_126 vdd gnd cell_6t
Xbit_r127_c146 bl_146 br_146 wl_127 vdd gnd cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd cell_6t
Xbit_r1_c147 bl_147 br_147 wl_1 vdd gnd cell_6t
Xbit_r2_c147 bl_147 br_147 wl_2 vdd gnd cell_6t
Xbit_r3_c147 bl_147 br_147 wl_3 vdd gnd cell_6t
Xbit_r4_c147 bl_147 br_147 wl_4 vdd gnd cell_6t
Xbit_r5_c147 bl_147 br_147 wl_5 vdd gnd cell_6t
Xbit_r6_c147 bl_147 br_147 wl_6 vdd gnd cell_6t
Xbit_r7_c147 bl_147 br_147 wl_7 vdd gnd cell_6t
Xbit_r8_c147 bl_147 br_147 wl_8 vdd gnd cell_6t
Xbit_r9_c147 bl_147 br_147 wl_9 vdd gnd cell_6t
Xbit_r10_c147 bl_147 br_147 wl_10 vdd gnd cell_6t
Xbit_r11_c147 bl_147 br_147 wl_11 vdd gnd cell_6t
Xbit_r12_c147 bl_147 br_147 wl_12 vdd gnd cell_6t
Xbit_r13_c147 bl_147 br_147 wl_13 vdd gnd cell_6t
Xbit_r14_c147 bl_147 br_147 wl_14 vdd gnd cell_6t
Xbit_r15_c147 bl_147 br_147 wl_15 vdd gnd cell_6t
Xbit_r16_c147 bl_147 br_147 wl_16 vdd gnd cell_6t
Xbit_r17_c147 bl_147 br_147 wl_17 vdd gnd cell_6t
Xbit_r18_c147 bl_147 br_147 wl_18 vdd gnd cell_6t
Xbit_r19_c147 bl_147 br_147 wl_19 vdd gnd cell_6t
Xbit_r20_c147 bl_147 br_147 wl_20 vdd gnd cell_6t
Xbit_r21_c147 bl_147 br_147 wl_21 vdd gnd cell_6t
Xbit_r22_c147 bl_147 br_147 wl_22 vdd gnd cell_6t
Xbit_r23_c147 bl_147 br_147 wl_23 vdd gnd cell_6t
Xbit_r24_c147 bl_147 br_147 wl_24 vdd gnd cell_6t
Xbit_r25_c147 bl_147 br_147 wl_25 vdd gnd cell_6t
Xbit_r26_c147 bl_147 br_147 wl_26 vdd gnd cell_6t
Xbit_r27_c147 bl_147 br_147 wl_27 vdd gnd cell_6t
Xbit_r28_c147 bl_147 br_147 wl_28 vdd gnd cell_6t
Xbit_r29_c147 bl_147 br_147 wl_29 vdd gnd cell_6t
Xbit_r30_c147 bl_147 br_147 wl_30 vdd gnd cell_6t
Xbit_r31_c147 bl_147 br_147 wl_31 vdd gnd cell_6t
Xbit_r32_c147 bl_147 br_147 wl_32 vdd gnd cell_6t
Xbit_r33_c147 bl_147 br_147 wl_33 vdd gnd cell_6t
Xbit_r34_c147 bl_147 br_147 wl_34 vdd gnd cell_6t
Xbit_r35_c147 bl_147 br_147 wl_35 vdd gnd cell_6t
Xbit_r36_c147 bl_147 br_147 wl_36 vdd gnd cell_6t
Xbit_r37_c147 bl_147 br_147 wl_37 vdd gnd cell_6t
Xbit_r38_c147 bl_147 br_147 wl_38 vdd gnd cell_6t
Xbit_r39_c147 bl_147 br_147 wl_39 vdd gnd cell_6t
Xbit_r40_c147 bl_147 br_147 wl_40 vdd gnd cell_6t
Xbit_r41_c147 bl_147 br_147 wl_41 vdd gnd cell_6t
Xbit_r42_c147 bl_147 br_147 wl_42 vdd gnd cell_6t
Xbit_r43_c147 bl_147 br_147 wl_43 vdd gnd cell_6t
Xbit_r44_c147 bl_147 br_147 wl_44 vdd gnd cell_6t
Xbit_r45_c147 bl_147 br_147 wl_45 vdd gnd cell_6t
Xbit_r46_c147 bl_147 br_147 wl_46 vdd gnd cell_6t
Xbit_r47_c147 bl_147 br_147 wl_47 vdd gnd cell_6t
Xbit_r48_c147 bl_147 br_147 wl_48 vdd gnd cell_6t
Xbit_r49_c147 bl_147 br_147 wl_49 vdd gnd cell_6t
Xbit_r50_c147 bl_147 br_147 wl_50 vdd gnd cell_6t
Xbit_r51_c147 bl_147 br_147 wl_51 vdd gnd cell_6t
Xbit_r52_c147 bl_147 br_147 wl_52 vdd gnd cell_6t
Xbit_r53_c147 bl_147 br_147 wl_53 vdd gnd cell_6t
Xbit_r54_c147 bl_147 br_147 wl_54 vdd gnd cell_6t
Xbit_r55_c147 bl_147 br_147 wl_55 vdd gnd cell_6t
Xbit_r56_c147 bl_147 br_147 wl_56 vdd gnd cell_6t
Xbit_r57_c147 bl_147 br_147 wl_57 vdd gnd cell_6t
Xbit_r58_c147 bl_147 br_147 wl_58 vdd gnd cell_6t
Xbit_r59_c147 bl_147 br_147 wl_59 vdd gnd cell_6t
Xbit_r60_c147 bl_147 br_147 wl_60 vdd gnd cell_6t
Xbit_r61_c147 bl_147 br_147 wl_61 vdd gnd cell_6t
Xbit_r62_c147 bl_147 br_147 wl_62 vdd gnd cell_6t
Xbit_r63_c147 bl_147 br_147 wl_63 vdd gnd cell_6t
Xbit_r64_c147 bl_147 br_147 wl_64 vdd gnd cell_6t
Xbit_r65_c147 bl_147 br_147 wl_65 vdd gnd cell_6t
Xbit_r66_c147 bl_147 br_147 wl_66 vdd gnd cell_6t
Xbit_r67_c147 bl_147 br_147 wl_67 vdd gnd cell_6t
Xbit_r68_c147 bl_147 br_147 wl_68 vdd gnd cell_6t
Xbit_r69_c147 bl_147 br_147 wl_69 vdd gnd cell_6t
Xbit_r70_c147 bl_147 br_147 wl_70 vdd gnd cell_6t
Xbit_r71_c147 bl_147 br_147 wl_71 vdd gnd cell_6t
Xbit_r72_c147 bl_147 br_147 wl_72 vdd gnd cell_6t
Xbit_r73_c147 bl_147 br_147 wl_73 vdd gnd cell_6t
Xbit_r74_c147 bl_147 br_147 wl_74 vdd gnd cell_6t
Xbit_r75_c147 bl_147 br_147 wl_75 vdd gnd cell_6t
Xbit_r76_c147 bl_147 br_147 wl_76 vdd gnd cell_6t
Xbit_r77_c147 bl_147 br_147 wl_77 vdd gnd cell_6t
Xbit_r78_c147 bl_147 br_147 wl_78 vdd gnd cell_6t
Xbit_r79_c147 bl_147 br_147 wl_79 vdd gnd cell_6t
Xbit_r80_c147 bl_147 br_147 wl_80 vdd gnd cell_6t
Xbit_r81_c147 bl_147 br_147 wl_81 vdd gnd cell_6t
Xbit_r82_c147 bl_147 br_147 wl_82 vdd gnd cell_6t
Xbit_r83_c147 bl_147 br_147 wl_83 vdd gnd cell_6t
Xbit_r84_c147 bl_147 br_147 wl_84 vdd gnd cell_6t
Xbit_r85_c147 bl_147 br_147 wl_85 vdd gnd cell_6t
Xbit_r86_c147 bl_147 br_147 wl_86 vdd gnd cell_6t
Xbit_r87_c147 bl_147 br_147 wl_87 vdd gnd cell_6t
Xbit_r88_c147 bl_147 br_147 wl_88 vdd gnd cell_6t
Xbit_r89_c147 bl_147 br_147 wl_89 vdd gnd cell_6t
Xbit_r90_c147 bl_147 br_147 wl_90 vdd gnd cell_6t
Xbit_r91_c147 bl_147 br_147 wl_91 vdd gnd cell_6t
Xbit_r92_c147 bl_147 br_147 wl_92 vdd gnd cell_6t
Xbit_r93_c147 bl_147 br_147 wl_93 vdd gnd cell_6t
Xbit_r94_c147 bl_147 br_147 wl_94 vdd gnd cell_6t
Xbit_r95_c147 bl_147 br_147 wl_95 vdd gnd cell_6t
Xbit_r96_c147 bl_147 br_147 wl_96 vdd gnd cell_6t
Xbit_r97_c147 bl_147 br_147 wl_97 vdd gnd cell_6t
Xbit_r98_c147 bl_147 br_147 wl_98 vdd gnd cell_6t
Xbit_r99_c147 bl_147 br_147 wl_99 vdd gnd cell_6t
Xbit_r100_c147 bl_147 br_147 wl_100 vdd gnd cell_6t
Xbit_r101_c147 bl_147 br_147 wl_101 vdd gnd cell_6t
Xbit_r102_c147 bl_147 br_147 wl_102 vdd gnd cell_6t
Xbit_r103_c147 bl_147 br_147 wl_103 vdd gnd cell_6t
Xbit_r104_c147 bl_147 br_147 wl_104 vdd gnd cell_6t
Xbit_r105_c147 bl_147 br_147 wl_105 vdd gnd cell_6t
Xbit_r106_c147 bl_147 br_147 wl_106 vdd gnd cell_6t
Xbit_r107_c147 bl_147 br_147 wl_107 vdd gnd cell_6t
Xbit_r108_c147 bl_147 br_147 wl_108 vdd gnd cell_6t
Xbit_r109_c147 bl_147 br_147 wl_109 vdd gnd cell_6t
Xbit_r110_c147 bl_147 br_147 wl_110 vdd gnd cell_6t
Xbit_r111_c147 bl_147 br_147 wl_111 vdd gnd cell_6t
Xbit_r112_c147 bl_147 br_147 wl_112 vdd gnd cell_6t
Xbit_r113_c147 bl_147 br_147 wl_113 vdd gnd cell_6t
Xbit_r114_c147 bl_147 br_147 wl_114 vdd gnd cell_6t
Xbit_r115_c147 bl_147 br_147 wl_115 vdd gnd cell_6t
Xbit_r116_c147 bl_147 br_147 wl_116 vdd gnd cell_6t
Xbit_r117_c147 bl_147 br_147 wl_117 vdd gnd cell_6t
Xbit_r118_c147 bl_147 br_147 wl_118 vdd gnd cell_6t
Xbit_r119_c147 bl_147 br_147 wl_119 vdd gnd cell_6t
Xbit_r120_c147 bl_147 br_147 wl_120 vdd gnd cell_6t
Xbit_r121_c147 bl_147 br_147 wl_121 vdd gnd cell_6t
Xbit_r122_c147 bl_147 br_147 wl_122 vdd gnd cell_6t
Xbit_r123_c147 bl_147 br_147 wl_123 vdd gnd cell_6t
Xbit_r124_c147 bl_147 br_147 wl_124 vdd gnd cell_6t
Xbit_r125_c147 bl_147 br_147 wl_125 vdd gnd cell_6t
Xbit_r126_c147 bl_147 br_147 wl_126 vdd gnd cell_6t
Xbit_r127_c147 bl_147 br_147 wl_127 vdd gnd cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd cell_6t
Xbit_r1_c148 bl_148 br_148 wl_1 vdd gnd cell_6t
Xbit_r2_c148 bl_148 br_148 wl_2 vdd gnd cell_6t
Xbit_r3_c148 bl_148 br_148 wl_3 vdd gnd cell_6t
Xbit_r4_c148 bl_148 br_148 wl_4 vdd gnd cell_6t
Xbit_r5_c148 bl_148 br_148 wl_5 vdd gnd cell_6t
Xbit_r6_c148 bl_148 br_148 wl_6 vdd gnd cell_6t
Xbit_r7_c148 bl_148 br_148 wl_7 vdd gnd cell_6t
Xbit_r8_c148 bl_148 br_148 wl_8 vdd gnd cell_6t
Xbit_r9_c148 bl_148 br_148 wl_9 vdd gnd cell_6t
Xbit_r10_c148 bl_148 br_148 wl_10 vdd gnd cell_6t
Xbit_r11_c148 bl_148 br_148 wl_11 vdd gnd cell_6t
Xbit_r12_c148 bl_148 br_148 wl_12 vdd gnd cell_6t
Xbit_r13_c148 bl_148 br_148 wl_13 vdd gnd cell_6t
Xbit_r14_c148 bl_148 br_148 wl_14 vdd gnd cell_6t
Xbit_r15_c148 bl_148 br_148 wl_15 vdd gnd cell_6t
Xbit_r16_c148 bl_148 br_148 wl_16 vdd gnd cell_6t
Xbit_r17_c148 bl_148 br_148 wl_17 vdd gnd cell_6t
Xbit_r18_c148 bl_148 br_148 wl_18 vdd gnd cell_6t
Xbit_r19_c148 bl_148 br_148 wl_19 vdd gnd cell_6t
Xbit_r20_c148 bl_148 br_148 wl_20 vdd gnd cell_6t
Xbit_r21_c148 bl_148 br_148 wl_21 vdd gnd cell_6t
Xbit_r22_c148 bl_148 br_148 wl_22 vdd gnd cell_6t
Xbit_r23_c148 bl_148 br_148 wl_23 vdd gnd cell_6t
Xbit_r24_c148 bl_148 br_148 wl_24 vdd gnd cell_6t
Xbit_r25_c148 bl_148 br_148 wl_25 vdd gnd cell_6t
Xbit_r26_c148 bl_148 br_148 wl_26 vdd gnd cell_6t
Xbit_r27_c148 bl_148 br_148 wl_27 vdd gnd cell_6t
Xbit_r28_c148 bl_148 br_148 wl_28 vdd gnd cell_6t
Xbit_r29_c148 bl_148 br_148 wl_29 vdd gnd cell_6t
Xbit_r30_c148 bl_148 br_148 wl_30 vdd gnd cell_6t
Xbit_r31_c148 bl_148 br_148 wl_31 vdd gnd cell_6t
Xbit_r32_c148 bl_148 br_148 wl_32 vdd gnd cell_6t
Xbit_r33_c148 bl_148 br_148 wl_33 vdd gnd cell_6t
Xbit_r34_c148 bl_148 br_148 wl_34 vdd gnd cell_6t
Xbit_r35_c148 bl_148 br_148 wl_35 vdd gnd cell_6t
Xbit_r36_c148 bl_148 br_148 wl_36 vdd gnd cell_6t
Xbit_r37_c148 bl_148 br_148 wl_37 vdd gnd cell_6t
Xbit_r38_c148 bl_148 br_148 wl_38 vdd gnd cell_6t
Xbit_r39_c148 bl_148 br_148 wl_39 vdd gnd cell_6t
Xbit_r40_c148 bl_148 br_148 wl_40 vdd gnd cell_6t
Xbit_r41_c148 bl_148 br_148 wl_41 vdd gnd cell_6t
Xbit_r42_c148 bl_148 br_148 wl_42 vdd gnd cell_6t
Xbit_r43_c148 bl_148 br_148 wl_43 vdd gnd cell_6t
Xbit_r44_c148 bl_148 br_148 wl_44 vdd gnd cell_6t
Xbit_r45_c148 bl_148 br_148 wl_45 vdd gnd cell_6t
Xbit_r46_c148 bl_148 br_148 wl_46 vdd gnd cell_6t
Xbit_r47_c148 bl_148 br_148 wl_47 vdd gnd cell_6t
Xbit_r48_c148 bl_148 br_148 wl_48 vdd gnd cell_6t
Xbit_r49_c148 bl_148 br_148 wl_49 vdd gnd cell_6t
Xbit_r50_c148 bl_148 br_148 wl_50 vdd gnd cell_6t
Xbit_r51_c148 bl_148 br_148 wl_51 vdd gnd cell_6t
Xbit_r52_c148 bl_148 br_148 wl_52 vdd gnd cell_6t
Xbit_r53_c148 bl_148 br_148 wl_53 vdd gnd cell_6t
Xbit_r54_c148 bl_148 br_148 wl_54 vdd gnd cell_6t
Xbit_r55_c148 bl_148 br_148 wl_55 vdd gnd cell_6t
Xbit_r56_c148 bl_148 br_148 wl_56 vdd gnd cell_6t
Xbit_r57_c148 bl_148 br_148 wl_57 vdd gnd cell_6t
Xbit_r58_c148 bl_148 br_148 wl_58 vdd gnd cell_6t
Xbit_r59_c148 bl_148 br_148 wl_59 vdd gnd cell_6t
Xbit_r60_c148 bl_148 br_148 wl_60 vdd gnd cell_6t
Xbit_r61_c148 bl_148 br_148 wl_61 vdd gnd cell_6t
Xbit_r62_c148 bl_148 br_148 wl_62 vdd gnd cell_6t
Xbit_r63_c148 bl_148 br_148 wl_63 vdd gnd cell_6t
Xbit_r64_c148 bl_148 br_148 wl_64 vdd gnd cell_6t
Xbit_r65_c148 bl_148 br_148 wl_65 vdd gnd cell_6t
Xbit_r66_c148 bl_148 br_148 wl_66 vdd gnd cell_6t
Xbit_r67_c148 bl_148 br_148 wl_67 vdd gnd cell_6t
Xbit_r68_c148 bl_148 br_148 wl_68 vdd gnd cell_6t
Xbit_r69_c148 bl_148 br_148 wl_69 vdd gnd cell_6t
Xbit_r70_c148 bl_148 br_148 wl_70 vdd gnd cell_6t
Xbit_r71_c148 bl_148 br_148 wl_71 vdd gnd cell_6t
Xbit_r72_c148 bl_148 br_148 wl_72 vdd gnd cell_6t
Xbit_r73_c148 bl_148 br_148 wl_73 vdd gnd cell_6t
Xbit_r74_c148 bl_148 br_148 wl_74 vdd gnd cell_6t
Xbit_r75_c148 bl_148 br_148 wl_75 vdd gnd cell_6t
Xbit_r76_c148 bl_148 br_148 wl_76 vdd gnd cell_6t
Xbit_r77_c148 bl_148 br_148 wl_77 vdd gnd cell_6t
Xbit_r78_c148 bl_148 br_148 wl_78 vdd gnd cell_6t
Xbit_r79_c148 bl_148 br_148 wl_79 vdd gnd cell_6t
Xbit_r80_c148 bl_148 br_148 wl_80 vdd gnd cell_6t
Xbit_r81_c148 bl_148 br_148 wl_81 vdd gnd cell_6t
Xbit_r82_c148 bl_148 br_148 wl_82 vdd gnd cell_6t
Xbit_r83_c148 bl_148 br_148 wl_83 vdd gnd cell_6t
Xbit_r84_c148 bl_148 br_148 wl_84 vdd gnd cell_6t
Xbit_r85_c148 bl_148 br_148 wl_85 vdd gnd cell_6t
Xbit_r86_c148 bl_148 br_148 wl_86 vdd gnd cell_6t
Xbit_r87_c148 bl_148 br_148 wl_87 vdd gnd cell_6t
Xbit_r88_c148 bl_148 br_148 wl_88 vdd gnd cell_6t
Xbit_r89_c148 bl_148 br_148 wl_89 vdd gnd cell_6t
Xbit_r90_c148 bl_148 br_148 wl_90 vdd gnd cell_6t
Xbit_r91_c148 bl_148 br_148 wl_91 vdd gnd cell_6t
Xbit_r92_c148 bl_148 br_148 wl_92 vdd gnd cell_6t
Xbit_r93_c148 bl_148 br_148 wl_93 vdd gnd cell_6t
Xbit_r94_c148 bl_148 br_148 wl_94 vdd gnd cell_6t
Xbit_r95_c148 bl_148 br_148 wl_95 vdd gnd cell_6t
Xbit_r96_c148 bl_148 br_148 wl_96 vdd gnd cell_6t
Xbit_r97_c148 bl_148 br_148 wl_97 vdd gnd cell_6t
Xbit_r98_c148 bl_148 br_148 wl_98 vdd gnd cell_6t
Xbit_r99_c148 bl_148 br_148 wl_99 vdd gnd cell_6t
Xbit_r100_c148 bl_148 br_148 wl_100 vdd gnd cell_6t
Xbit_r101_c148 bl_148 br_148 wl_101 vdd gnd cell_6t
Xbit_r102_c148 bl_148 br_148 wl_102 vdd gnd cell_6t
Xbit_r103_c148 bl_148 br_148 wl_103 vdd gnd cell_6t
Xbit_r104_c148 bl_148 br_148 wl_104 vdd gnd cell_6t
Xbit_r105_c148 bl_148 br_148 wl_105 vdd gnd cell_6t
Xbit_r106_c148 bl_148 br_148 wl_106 vdd gnd cell_6t
Xbit_r107_c148 bl_148 br_148 wl_107 vdd gnd cell_6t
Xbit_r108_c148 bl_148 br_148 wl_108 vdd gnd cell_6t
Xbit_r109_c148 bl_148 br_148 wl_109 vdd gnd cell_6t
Xbit_r110_c148 bl_148 br_148 wl_110 vdd gnd cell_6t
Xbit_r111_c148 bl_148 br_148 wl_111 vdd gnd cell_6t
Xbit_r112_c148 bl_148 br_148 wl_112 vdd gnd cell_6t
Xbit_r113_c148 bl_148 br_148 wl_113 vdd gnd cell_6t
Xbit_r114_c148 bl_148 br_148 wl_114 vdd gnd cell_6t
Xbit_r115_c148 bl_148 br_148 wl_115 vdd gnd cell_6t
Xbit_r116_c148 bl_148 br_148 wl_116 vdd gnd cell_6t
Xbit_r117_c148 bl_148 br_148 wl_117 vdd gnd cell_6t
Xbit_r118_c148 bl_148 br_148 wl_118 vdd gnd cell_6t
Xbit_r119_c148 bl_148 br_148 wl_119 vdd gnd cell_6t
Xbit_r120_c148 bl_148 br_148 wl_120 vdd gnd cell_6t
Xbit_r121_c148 bl_148 br_148 wl_121 vdd gnd cell_6t
Xbit_r122_c148 bl_148 br_148 wl_122 vdd gnd cell_6t
Xbit_r123_c148 bl_148 br_148 wl_123 vdd gnd cell_6t
Xbit_r124_c148 bl_148 br_148 wl_124 vdd gnd cell_6t
Xbit_r125_c148 bl_148 br_148 wl_125 vdd gnd cell_6t
Xbit_r126_c148 bl_148 br_148 wl_126 vdd gnd cell_6t
Xbit_r127_c148 bl_148 br_148 wl_127 vdd gnd cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd cell_6t
Xbit_r1_c149 bl_149 br_149 wl_1 vdd gnd cell_6t
Xbit_r2_c149 bl_149 br_149 wl_2 vdd gnd cell_6t
Xbit_r3_c149 bl_149 br_149 wl_3 vdd gnd cell_6t
Xbit_r4_c149 bl_149 br_149 wl_4 vdd gnd cell_6t
Xbit_r5_c149 bl_149 br_149 wl_5 vdd gnd cell_6t
Xbit_r6_c149 bl_149 br_149 wl_6 vdd gnd cell_6t
Xbit_r7_c149 bl_149 br_149 wl_7 vdd gnd cell_6t
Xbit_r8_c149 bl_149 br_149 wl_8 vdd gnd cell_6t
Xbit_r9_c149 bl_149 br_149 wl_9 vdd gnd cell_6t
Xbit_r10_c149 bl_149 br_149 wl_10 vdd gnd cell_6t
Xbit_r11_c149 bl_149 br_149 wl_11 vdd gnd cell_6t
Xbit_r12_c149 bl_149 br_149 wl_12 vdd gnd cell_6t
Xbit_r13_c149 bl_149 br_149 wl_13 vdd gnd cell_6t
Xbit_r14_c149 bl_149 br_149 wl_14 vdd gnd cell_6t
Xbit_r15_c149 bl_149 br_149 wl_15 vdd gnd cell_6t
Xbit_r16_c149 bl_149 br_149 wl_16 vdd gnd cell_6t
Xbit_r17_c149 bl_149 br_149 wl_17 vdd gnd cell_6t
Xbit_r18_c149 bl_149 br_149 wl_18 vdd gnd cell_6t
Xbit_r19_c149 bl_149 br_149 wl_19 vdd gnd cell_6t
Xbit_r20_c149 bl_149 br_149 wl_20 vdd gnd cell_6t
Xbit_r21_c149 bl_149 br_149 wl_21 vdd gnd cell_6t
Xbit_r22_c149 bl_149 br_149 wl_22 vdd gnd cell_6t
Xbit_r23_c149 bl_149 br_149 wl_23 vdd gnd cell_6t
Xbit_r24_c149 bl_149 br_149 wl_24 vdd gnd cell_6t
Xbit_r25_c149 bl_149 br_149 wl_25 vdd gnd cell_6t
Xbit_r26_c149 bl_149 br_149 wl_26 vdd gnd cell_6t
Xbit_r27_c149 bl_149 br_149 wl_27 vdd gnd cell_6t
Xbit_r28_c149 bl_149 br_149 wl_28 vdd gnd cell_6t
Xbit_r29_c149 bl_149 br_149 wl_29 vdd gnd cell_6t
Xbit_r30_c149 bl_149 br_149 wl_30 vdd gnd cell_6t
Xbit_r31_c149 bl_149 br_149 wl_31 vdd gnd cell_6t
Xbit_r32_c149 bl_149 br_149 wl_32 vdd gnd cell_6t
Xbit_r33_c149 bl_149 br_149 wl_33 vdd gnd cell_6t
Xbit_r34_c149 bl_149 br_149 wl_34 vdd gnd cell_6t
Xbit_r35_c149 bl_149 br_149 wl_35 vdd gnd cell_6t
Xbit_r36_c149 bl_149 br_149 wl_36 vdd gnd cell_6t
Xbit_r37_c149 bl_149 br_149 wl_37 vdd gnd cell_6t
Xbit_r38_c149 bl_149 br_149 wl_38 vdd gnd cell_6t
Xbit_r39_c149 bl_149 br_149 wl_39 vdd gnd cell_6t
Xbit_r40_c149 bl_149 br_149 wl_40 vdd gnd cell_6t
Xbit_r41_c149 bl_149 br_149 wl_41 vdd gnd cell_6t
Xbit_r42_c149 bl_149 br_149 wl_42 vdd gnd cell_6t
Xbit_r43_c149 bl_149 br_149 wl_43 vdd gnd cell_6t
Xbit_r44_c149 bl_149 br_149 wl_44 vdd gnd cell_6t
Xbit_r45_c149 bl_149 br_149 wl_45 vdd gnd cell_6t
Xbit_r46_c149 bl_149 br_149 wl_46 vdd gnd cell_6t
Xbit_r47_c149 bl_149 br_149 wl_47 vdd gnd cell_6t
Xbit_r48_c149 bl_149 br_149 wl_48 vdd gnd cell_6t
Xbit_r49_c149 bl_149 br_149 wl_49 vdd gnd cell_6t
Xbit_r50_c149 bl_149 br_149 wl_50 vdd gnd cell_6t
Xbit_r51_c149 bl_149 br_149 wl_51 vdd gnd cell_6t
Xbit_r52_c149 bl_149 br_149 wl_52 vdd gnd cell_6t
Xbit_r53_c149 bl_149 br_149 wl_53 vdd gnd cell_6t
Xbit_r54_c149 bl_149 br_149 wl_54 vdd gnd cell_6t
Xbit_r55_c149 bl_149 br_149 wl_55 vdd gnd cell_6t
Xbit_r56_c149 bl_149 br_149 wl_56 vdd gnd cell_6t
Xbit_r57_c149 bl_149 br_149 wl_57 vdd gnd cell_6t
Xbit_r58_c149 bl_149 br_149 wl_58 vdd gnd cell_6t
Xbit_r59_c149 bl_149 br_149 wl_59 vdd gnd cell_6t
Xbit_r60_c149 bl_149 br_149 wl_60 vdd gnd cell_6t
Xbit_r61_c149 bl_149 br_149 wl_61 vdd gnd cell_6t
Xbit_r62_c149 bl_149 br_149 wl_62 vdd gnd cell_6t
Xbit_r63_c149 bl_149 br_149 wl_63 vdd gnd cell_6t
Xbit_r64_c149 bl_149 br_149 wl_64 vdd gnd cell_6t
Xbit_r65_c149 bl_149 br_149 wl_65 vdd gnd cell_6t
Xbit_r66_c149 bl_149 br_149 wl_66 vdd gnd cell_6t
Xbit_r67_c149 bl_149 br_149 wl_67 vdd gnd cell_6t
Xbit_r68_c149 bl_149 br_149 wl_68 vdd gnd cell_6t
Xbit_r69_c149 bl_149 br_149 wl_69 vdd gnd cell_6t
Xbit_r70_c149 bl_149 br_149 wl_70 vdd gnd cell_6t
Xbit_r71_c149 bl_149 br_149 wl_71 vdd gnd cell_6t
Xbit_r72_c149 bl_149 br_149 wl_72 vdd gnd cell_6t
Xbit_r73_c149 bl_149 br_149 wl_73 vdd gnd cell_6t
Xbit_r74_c149 bl_149 br_149 wl_74 vdd gnd cell_6t
Xbit_r75_c149 bl_149 br_149 wl_75 vdd gnd cell_6t
Xbit_r76_c149 bl_149 br_149 wl_76 vdd gnd cell_6t
Xbit_r77_c149 bl_149 br_149 wl_77 vdd gnd cell_6t
Xbit_r78_c149 bl_149 br_149 wl_78 vdd gnd cell_6t
Xbit_r79_c149 bl_149 br_149 wl_79 vdd gnd cell_6t
Xbit_r80_c149 bl_149 br_149 wl_80 vdd gnd cell_6t
Xbit_r81_c149 bl_149 br_149 wl_81 vdd gnd cell_6t
Xbit_r82_c149 bl_149 br_149 wl_82 vdd gnd cell_6t
Xbit_r83_c149 bl_149 br_149 wl_83 vdd gnd cell_6t
Xbit_r84_c149 bl_149 br_149 wl_84 vdd gnd cell_6t
Xbit_r85_c149 bl_149 br_149 wl_85 vdd gnd cell_6t
Xbit_r86_c149 bl_149 br_149 wl_86 vdd gnd cell_6t
Xbit_r87_c149 bl_149 br_149 wl_87 vdd gnd cell_6t
Xbit_r88_c149 bl_149 br_149 wl_88 vdd gnd cell_6t
Xbit_r89_c149 bl_149 br_149 wl_89 vdd gnd cell_6t
Xbit_r90_c149 bl_149 br_149 wl_90 vdd gnd cell_6t
Xbit_r91_c149 bl_149 br_149 wl_91 vdd gnd cell_6t
Xbit_r92_c149 bl_149 br_149 wl_92 vdd gnd cell_6t
Xbit_r93_c149 bl_149 br_149 wl_93 vdd gnd cell_6t
Xbit_r94_c149 bl_149 br_149 wl_94 vdd gnd cell_6t
Xbit_r95_c149 bl_149 br_149 wl_95 vdd gnd cell_6t
Xbit_r96_c149 bl_149 br_149 wl_96 vdd gnd cell_6t
Xbit_r97_c149 bl_149 br_149 wl_97 vdd gnd cell_6t
Xbit_r98_c149 bl_149 br_149 wl_98 vdd gnd cell_6t
Xbit_r99_c149 bl_149 br_149 wl_99 vdd gnd cell_6t
Xbit_r100_c149 bl_149 br_149 wl_100 vdd gnd cell_6t
Xbit_r101_c149 bl_149 br_149 wl_101 vdd gnd cell_6t
Xbit_r102_c149 bl_149 br_149 wl_102 vdd gnd cell_6t
Xbit_r103_c149 bl_149 br_149 wl_103 vdd gnd cell_6t
Xbit_r104_c149 bl_149 br_149 wl_104 vdd gnd cell_6t
Xbit_r105_c149 bl_149 br_149 wl_105 vdd gnd cell_6t
Xbit_r106_c149 bl_149 br_149 wl_106 vdd gnd cell_6t
Xbit_r107_c149 bl_149 br_149 wl_107 vdd gnd cell_6t
Xbit_r108_c149 bl_149 br_149 wl_108 vdd gnd cell_6t
Xbit_r109_c149 bl_149 br_149 wl_109 vdd gnd cell_6t
Xbit_r110_c149 bl_149 br_149 wl_110 vdd gnd cell_6t
Xbit_r111_c149 bl_149 br_149 wl_111 vdd gnd cell_6t
Xbit_r112_c149 bl_149 br_149 wl_112 vdd gnd cell_6t
Xbit_r113_c149 bl_149 br_149 wl_113 vdd gnd cell_6t
Xbit_r114_c149 bl_149 br_149 wl_114 vdd gnd cell_6t
Xbit_r115_c149 bl_149 br_149 wl_115 vdd gnd cell_6t
Xbit_r116_c149 bl_149 br_149 wl_116 vdd gnd cell_6t
Xbit_r117_c149 bl_149 br_149 wl_117 vdd gnd cell_6t
Xbit_r118_c149 bl_149 br_149 wl_118 vdd gnd cell_6t
Xbit_r119_c149 bl_149 br_149 wl_119 vdd gnd cell_6t
Xbit_r120_c149 bl_149 br_149 wl_120 vdd gnd cell_6t
Xbit_r121_c149 bl_149 br_149 wl_121 vdd gnd cell_6t
Xbit_r122_c149 bl_149 br_149 wl_122 vdd gnd cell_6t
Xbit_r123_c149 bl_149 br_149 wl_123 vdd gnd cell_6t
Xbit_r124_c149 bl_149 br_149 wl_124 vdd gnd cell_6t
Xbit_r125_c149 bl_149 br_149 wl_125 vdd gnd cell_6t
Xbit_r126_c149 bl_149 br_149 wl_126 vdd gnd cell_6t
Xbit_r127_c149 bl_149 br_149 wl_127 vdd gnd cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd cell_6t
Xbit_r1_c150 bl_150 br_150 wl_1 vdd gnd cell_6t
Xbit_r2_c150 bl_150 br_150 wl_2 vdd gnd cell_6t
Xbit_r3_c150 bl_150 br_150 wl_3 vdd gnd cell_6t
Xbit_r4_c150 bl_150 br_150 wl_4 vdd gnd cell_6t
Xbit_r5_c150 bl_150 br_150 wl_5 vdd gnd cell_6t
Xbit_r6_c150 bl_150 br_150 wl_6 vdd gnd cell_6t
Xbit_r7_c150 bl_150 br_150 wl_7 vdd gnd cell_6t
Xbit_r8_c150 bl_150 br_150 wl_8 vdd gnd cell_6t
Xbit_r9_c150 bl_150 br_150 wl_9 vdd gnd cell_6t
Xbit_r10_c150 bl_150 br_150 wl_10 vdd gnd cell_6t
Xbit_r11_c150 bl_150 br_150 wl_11 vdd gnd cell_6t
Xbit_r12_c150 bl_150 br_150 wl_12 vdd gnd cell_6t
Xbit_r13_c150 bl_150 br_150 wl_13 vdd gnd cell_6t
Xbit_r14_c150 bl_150 br_150 wl_14 vdd gnd cell_6t
Xbit_r15_c150 bl_150 br_150 wl_15 vdd gnd cell_6t
Xbit_r16_c150 bl_150 br_150 wl_16 vdd gnd cell_6t
Xbit_r17_c150 bl_150 br_150 wl_17 vdd gnd cell_6t
Xbit_r18_c150 bl_150 br_150 wl_18 vdd gnd cell_6t
Xbit_r19_c150 bl_150 br_150 wl_19 vdd gnd cell_6t
Xbit_r20_c150 bl_150 br_150 wl_20 vdd gnd cell_6t
Xbit_r21_c150 bl_150 br_150 wl_21 vdd gnd cell_6t
Xbit_r22_c150 bl_150 br_150 wl_22 vdd gnd cell_6t
Xbit_r23_c150 bl_150 br_150 wl_23 vdd gnd cell_6t
Xbit_r24_c150 bl_150 br_150 wl_24 vdd gnd cell_6t
Xbit_r25_c150 bl_150 br_150 wl_25 vdd gnd cell_6t
Xbit_r26_c150 bl_150 br_150 wl_26 vdd gnd cell_6t
Xbit_r27_c150 bl_150 br_150 wl_27 vdd gnd cell_6t
Xbit_r28_c150 bl_150 br_150 wl_28 vdd gnd cell_6t
Xbit_r29_c150 bl_150 br_150 wl_29 vdd gnd cell_6t
Xbit_r30_c150 bl_150 br_150 wl_30 vdd gnd cell_6t
Xbit_r31_c150 bl_150 br_150 wl_31 vdd gnd cell_6t
Xbit_r32_c150 bl_150 br_150 wl_32 vdd gnd cell_6t
Xbit_r33_c150 bl_150 br_150 wl_33 vdd gnd cell_6t
Xbit_r34_c150 bl_150 br_150 wl_34 vdd gnd cell_6t
Xbit_r35_c150 bl_150 br_150 wl_35 vdd gnd cell_6t
Xbit_r36_c150 bl_150 br_150 wl_36 vdd gnd cell_6t
Xbit_r37_c150 bl_150 br_150 wl_37 vdd gnd cell_6t
Xbit_r38_c150 bl_150 br_150 wl_38 vdd gnd cell_6t
Xbit_r39_c150 bl_150 br_150 wl_39 vdd gnd cell_6t
Xbit_r40_c150 bl_150 br_150 wl_40 vdd gnd cell_6t
Xbit_r41_c150 bl_150 br_150 wl_41 vdd gnd cell_6t
Xbit_r42_c150 bl_150 br_150 wl_42 vdd gnd cell_6t
Xbit_r43_c150 bl_150 br_150 wl_43 vdd gnd cell_6t
Xbit_r44_c150 bl_150 br_150 wl_44 vdd gnd cell_6t
Xbit_r45_c150 bl_150 br_150 wl_45 vdd gnd cell_6t
Xbit_r46_c150 bl_150 br_150 wl_46 vdd gnd cell_6t
Xbit_r47_c150 bl_150 br_150 wl_47 vdd gnd cell_6t
Xbit_r48_c150 bl_150 br_150 wl_48 vdd gnd cell_6t
Xbit_r49_c150 bl_150 br_150 wl_49 vdd gnd cell_6t
Xbit_r50_c150 bl_150 br_150 wl_50 vdd gnd cell_6t
Xbit_r51_c150 bl_150 br_150 wl_51 vdd gnd cell_6t
Xbit_r52_c150 bl_150 br_150 wl_52 vdd gnd cell_6t
Xbit_r53_c150 bl_150 br_150 wl_53 vdd gnd cell_6t
Xbit_r54_c150 bl_150 br_150 wl_54 vdd gnd cell_6t
Xbit_r55_c150 bl_150 br_150 wl_55 vdd gnd cell_6t
Xbit_r56_c150 bl_150 br_150 wl_56 vdd gnd cell_6t
Xbit_r57_c150 bl_150 br_150 wl_57 vdd gnd cell_6t
Xbit_r58_c150 bl_150 br_150 wl_58 vdd gnd cell_6t
Xbit_r59_c150 bl_150 br_150 wl_59 vdd gnd cell_6t
Xbit_r60_c150 bl_150 br_150 wl_60 vdd gnd cell_6t
Xbit_r61_c150 bl_150 br_150 wl_61 vdd gnd cell_6t
Xbit_r62_c150 bl_150 br_150 wl_62 vdd gnd cell_6t
Xbit_r63_c150 bl_150 br_150 wl_63 vdd gnd cell_6t
Xbit_r64_c150 bl_150 br_150 wl_64 vdd gnd cell_6t
Xbit_r65_c150 bl_150 br_150 wl_65 vdd gnd cell_6t
Xbit_r66_c150 bl_150 br_150 wl_66 vdd gnd cell_6t
Xbit_r67_c150 bl_150 br_150 wl_67 vdd gnd cell_6t
Xbit_r68_c150 bl_150 br_150 wl_68 vdd gnd cell_6t
Xbit_r69_c150 bl_150 br_150 wl_69 vdd gnd cell_6t
Xbit_r70_c150 bl_150 br_150 wl_70 vdd gnd cell_6t
Xbit_r71_c150 bl_150 br_150 wl_71 vdd gnd cell_6t
Xbit_r72_c150 bl_150 br_150 wl_72 vdd gnd cell_6t
Xbit_r73_c150 bl_150 br_150 wl_73 vdd gnd cell_6t
Xbit_r74_c150 bl_150 br_150 wl_74 vdd gnd cell_6t
Xbit_r75_c150 bl_150 br_150 wl_75 vdd gnd cell_6t
Xbit_r76_c150 bl_150 br_150 wl_76 vdd gnd cell_6t
Xbit_r77_c150 bl_150 br_150 wl_77 vdd gnd cell_6t
Xbit_r78_c150 bl_150 br_150 wl_78 vdd gnd cell_6t
Xbit_r79_c150 bl_150 br_150 wl_79 vdd gnd cell_6t
Xbit_r80_c150 bl_150 br_150 wl_80 vdd gnd cell_6t
Xbit_r81_c150 bl_150 br_150 wl_81 vdd gnd cell_6t
Xbit_r82_c150 bl_150 br_150 wl_82 vdd gnd cell_6t
Xbit_r83_c150 bl_150 br_150 wl_83 vdd gnd cell_6t
Xbit_r84_c150 bl_150 br_150 wl_84 vdd gnd cell_6t
Xbit_r85_c150 bl_150 br_150 wl_85 vdd gnd cell_6t
Xbit_r86_c150 bl_150 br_150 wl_86 vdd gnd cell_6t
Xbit_r87_c150 bl_150 br_150 wl_87 vdd gnd cell_6t
Xbit_r88_c150 bl_150 br_150 wl_88 vdd gnd cell_6t
Xbit_r89_c150 bl_150 br_150 wl_89 vdd gnd cell_6t
Xbit_r90_c150 bl_150 br_150 wl_90 vdd gnd cell_6t
Xbit_r91_c150 bl_150 br_150 wl_91 vdd gnd cell_6t
Xbit_r92_c150 bl_150 br_150 wl_92 vdd gnd cell_6t
Xbit_r93_c150 bl_150 br_150 wl_93 vdd gnd cell_6t
Xbit_r94_c150 bl_150 br_150 wl_94 vdd gnd cell_6t
Xbit_r95_c150 bl_150 br_150 wl_95 vdd gnd cell_6t
Xbit_r96_c150 bl_150 br_150 wl_96 vdd gnd cell_6t
Xbit_r97_c150 bl_150 br_150 wl_97 vdd gnd cell_6t
Xbit_r98_c150 bl_150 br_150 wl_98 vdd gnd cell_6t
Xbit_r99_c150 bl_150 br_150 wl_99 vdd gnd cell_6t
Xbit_r100_c150 bl_150 br_150 wl_100 vdd gnd cell_6t
Xbit_r101_c150 bl_150 br_150 wl_101 vdd gnd cell_6t
Xbit_r102_c150 bl_150 br_150 wl_102 vdd gnd cell_6t
Xbit_r103_c150 bl_150 br_150 wl_103 vdd gnd cell_6t
Xbit_r104_c150 bl_150 br_150 wl_104 vdd gnd cell_6t
Xbit_r105_c150 bl_150 br_150 wl_105 vdd gnd cell_6t
Xbit_r106_c150 bl_150 br_150 wl_106 vdd gnd cell_6t
Xbit_r107_c150 bl_150 br_150 wl_107 vdd gnd cell_6t
Xbit_r108_c150 bl_150 br_150 wl_108 vdd gnd cell_6t
Xbit_r109_c150 bl_150 br_150 wl_109 vdd gnd cell_6t
Xbit_r110_c150 bl_150 br_150 wl_110 vdd gnd cell_6t
Xbit_r111_c150 bl_150 br_150 wl_111 vdd gnd cell_6t
Xbit_r112_c150 bl_150 br_150 wl_112 vdd gnd cell_6t
Xbit_r113_c150 bl_150 br_150 wl_113 vdd gnd cell_6t
Xbit_r114_c150 bl_150 br_150 wl_114 vdd gnd cell_6t
Xbit_r115_c150 bl_150 br_150 wl_115 vdd gnd cell_6t
Xbit_r116_c150 bl_150 br_150 wl_116 vdd gnd cell_6t
Xbit_r117_c150 bl_150 br_150 wl_117 vdd gnd cell_6t
Xbit_r118_c150 bl_150 br_150 wl_118 vdd gnd cell_6t
Xbit_r119_c150 bl_150 br_150 wl_119 vdd gnd cell_6t
Xbit_r120_c150 bl_150 br_150 wl_120 vdd gnd cell_6t
Xbit_r121_c150 bl_150 br_150 wl_121 vdd gnd cell_6t
Xbit_r122_c150 bl_150 br_150 wl_122 vdd gnd cell_6t
Xbit_r123_c150 bl_150 br_150 wl_123 vdd gnd cell_6t
Xbit_r124_c150 bl_150 br_150 wl_124 vdd gnd cell_6t
Xbit_r125_c150 bl_150 br_150 wl_125 vdd gnd cell_6t
Xbit_r126_c150 bl_150 br_150 wl_126 vdd gnd cell_6t
Xbit_r127_c150 bl_150 br_150 wl_127 vdd gnd cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd cell_6t
Xbit_r1_c151 bl_151 br_151 wl_1 vdd gnd cell_6t
Xbit_r2_c151 bl_151 br_151 wl_2 vdd gnd cell_6t
Xbit_r3_c151 bl_151 br_151 wl_3 vdd gnd cell_6t
Xbit_r4_c151 bl_151 br_151 wl_4 vdd gnd cell_6t
Xbit_r5_c151 bl_151 br_151 wl_5 vdd gnd cell_6t
Xbit_r6_c151 bl_151 br_151 wl_6 vdd gnd cell_6t
Xbit_r7_c151 bl_151 br_151 wl_7 vdd gnd cell_6t
Xbit_r8_c151 bl_151 br_151 wl_8 vdd gnd cell_6t
Xbit_r9_c151 bl_151 br_151 wl_9 vdd gnd cell_6t
Xbit_r10_c151 bl_151 br_151 wl_10 vdd gnd cell_6t
Xbit_r11_c151 bl_151 br_151 wl_11 vdd gnd cell_6t
Xbit_r12_c151 bl_151 br_151 wl_12 vdd gnd cell_6t
Xbit_r13_c151 bl_151 br_151 wl_13 vdd gnd cell_6t
Xbit_r14_c151 bl_151 br_151 wl_14 vdd gnd cell_6t
Xbit_r15_c151 bl_151 br_151 wl_15 vdd gnd cell_6t
Xbit_r16_c151 bl_151 br_151 wl_16 vdd gnd cell_6t
Xbit_r17_c151 bl_151 br_151 wl_17 vdd gnd cell_6t
Xbit_r18_c151 bl_151 br_151 wl_18 vdd gnd cell_6t
Xbit_r19_c151 bl_151 br_151 wl_19 vdd gnd cell_6t
Xbit_r20_c151 bl_151 br_151 wl_20 vdd gnd cell_6t
Xbit_r21_c151 bl_151 br_151 wl_21 vdd gnd cell_6t
Xbit_r22_c151 bl_151 br_151 wl_22 vdd gnd cell_6t
Xbit_r23_c151 bl_151 br_151 wl_23 vdd gnd cell_6t
Xbit_r24_c151 bl_151 br_151 wl_24 vdd gnd cell_6t
Xbit_r25_c151 bl_151 br_151 wl_25 vdd gnd cell_6t
Xbit_r26_c151 bl_151 br_151 wl_26 vdd gnd cell_6t
Xbit_r27_c151 bl_151 br_151 wl_27 vdd gnd cell_6t
Xbit_r28_c151 bl_151 br_151 wl_28 vdd gnd cell_6t
Xbit_r29_c151 bl_151 br_151 wl_29 vdd gnd cell_6t
Xbit_r30_c151 bl_151 br_151 wl_30 vdd gnd cell_6t
Xbit_r31_c151 bl_151 br_151 wl_31 vdd gnd cell_6t
Xbit_r32_c151 bl_151 br_151 wl_32 vdd gnd cell_6t
Xbit_r33_c151 bl_151 br_151 wl_33 vdd gnd cell_6t
Xbit_r34_c151 bl_151 br_151 wl_34 vdd gnd cell_6t
Xbit_r35_c151 bl_151 br_151 wl_35 vdd gnd cell_6t
Xbit_r36_c151 bl_151 br_151 wl_36 vdd gnd cell_6t
Xbit_r37_c151 bl_151 br_151 wl_37 vdd gnd cell_6t
Xbit_r38_c151 bl_151 br_151 wl_38 vdd gnd cell_6t
Xbit_r39_c151 bl_151 br_151 wl_39 vdd gnd cell_6t
Xbit_r40_c151 bl_151 br_151 wl_40 vdd gnd cell_6t
Xbit_r41_c151 bl_151 br_151 wl_41 vdd gnd cell_6t
Xbit_r42_c151 bl_151 br_151 wl_42 vdd gnd cell_6t
Xbit_r43_c151 bl_151 br_151 wl_43 vdd gnd cell_6t
Xbit_r44_c151 bl_151 br_151 wl_44 vdd gnd cell_6t
Xbit_r45_c151 bl_151 br_151 wl_45 vdd gnd cell_6t
Xbit_r46_c151 bl_151 br_151 wl_46 vdd gnd cell_6t
Xbit_r47_c151 bl_151 br_151 wl_47 vdd gnd cell_6t
Xbit_r48_c151 bl_151 br_151 wl_48 vdd gnd cell_6t
Xbit_r49_c151 bl_151 br_151 wl_49 vdd gnd cell_6t
Xbit_r50_c151 bl_151 br_151 wl_50 vdd gnd cell_6t
Xbit_r51_c151 bl_151 br_151 wl_51 vdd gnd cell_6t
Xbit_r52_c151 bl_151 br_151 wl_52 vdd gnd cell_6t
Xbit_r53_c151 bl_151 br_151 wl_53 vdd gnd cell_6t
Xbit_r54_c151 bl_151 br_151 wl_54 vdd gnd cell_6t
Xbit_r55_c151 bl_151 br_151 wl_55 vdd gnd cell_6t
Xbit_r56_c151 bl_151 br_151 wl_56 vdd gnd cell_6t
Xbit_r57_c151 bl_151 br_151 wl_57 vdd gnd cell_6t
Xbit_r58_c151 bl_151 br_151 wl_58 vdd gnd cell_6t
Xbit_r59_c151 bl_151 br_151 wl_59 vdd gnd cell_6t
Xbit_r60_c151 bl_151 br_151 wl_60 vdd gnd cell_6t
Xbit_r61_c151 bl_151 br_151 wl_61 vdd gnd cell_6t
Xbit_r62_c151 bl_151 br_151 wl_62 vdd gnd cell_6t
Xbit_r63_c151 bl_151 br_151 wl_63 vdd gnd cell_6t
Xbit_r64_c151 bl_151 br_151 wl_64 vdd gnd cell_6t
Xbit_r65_c151 bl_151 br_151 wl_65 vdd gnd cell_6t
Xbit_r66_c151 bl_151 br_151 wl_66 vdd gnd cell_6t
Xbit_r67_c151 bl_151 br_151 wl_67 vdd gnd cell_6t
Xbit_r68_c151 bl_151 br_151 wl_68 vdd gnd cell_6t
Xbit_r69_c151 bl_151 br_151 wl_69 vdd gnd cell_6t
Xbit_r70_c151 bl_151 br_151 wl_70 vdd gnd cell_6t
Xbit_r71_c151 bl_151 br_151 wl_71 vdd gnd cell_6t
Xbit_r72_c151 bl_151 br_151 wl_72 vdd gnd cell_6t
Xbit_r73_c151 bl_151 br_151 wl_73 vdd gnd cell_6t
Xbit_r74_c151 bl_151 br_151 wl_74 vdd gnd cell_6t
Xbit_r75_c151 bl_151 br_151 wl_75 vdd gnd cell_6t
Xbit_r76_c151 bl_151 br_151 wl_76 vdd gnd cell_6t
Xbit_r77_c151 bl_151 br_151 wl_77 vdd gnd cell_6t
Xbit_r78_c151 bl_151 br_151 wl_78 vdd gnd cell_6t
Xbit_r79_c151 bl_151 br_151 wl_79 vdd gnd cell_6t
Xbit_r80_c151 bl_151 br_151 wl_80 vdd gnd cell_6t
Xbit_r81_c151 bl_151 br_151 wl_81 vdd gnd cell_6t
Xbit_r82_c151 bl_151 br_151 wl_82 vdd gnd cell_6t
Xbit_r83_c151 bl_151 br_151 wl_83 vdd gnd cell_6t
Xbit_r84_c151 bl_151 br_151 wl_84 vdd gnd cell_6t
Xbit_r85_c151 bl_151 br_151 wl_85 vdd gnd cell_6t
Xbit_r86_c151 bl_151 br_151 wl_86 vdd gnd cell_6t
Xbit_r87_c151 bl_151 br_151 wl_87 vdd gnd cell_6t
Xbit_r88_c151 bl_151 br_151 wl_88 vdd gnd cell_6t
Xbit_r89_c151 bl_151 br_151 wl_89 vdd gnd cell_6t
Xbit_r90_c151 bl_151 br_151 wl_90 vdd gnd cell_6t
Xbit_r91_c151 bl_151 br_151 wl_91 vdd gnd cell_6t
Xbit_r92_c151 bl_151 br_151 wl_92 vdd gnd cell_6t
Xbit_r93_c151 bl_151 br_151 wl_93 vdd gnd cell_6t
Xbit_r94_c151 bl_151 br_151 wl_94 vdd gnd cell_6t
Xbit_r95_c151 bl_151 br_151 wl_95 vdd gnd cell_6t
Xbit_r96_c151 bl_151 br_151 wl_96 vdd gnd cell_6t
Xbit_r97_c151 bl_151 br_151 wl_97 vdd gnd cell_6t
Xbit_r98_c151 bl_151 br_151 wl_98 vdd gnd cell_6t
Xbit_r99_c151 bl_151 br_151 wl_99 vdd gnd cell_6t
Xbit_r100_c151 bl_151 br_151 wl_100 vdd gnd cell_6t
Xbit_r101_c151 bl_151 br_151 wl_101 vdd gnd cell_6t
Xbit_r102_c151 bl_151 br_151 wl_102 vdd gnd cell_6t
Xbit_r103_c151 bl_151 br_151 wl_103 vdd gnd cell_6t
Xbit_r104_c151 bl_151 br_151 wl_104 vdd gnd cell_6t
Xbit_r105_c151 bl_151 br_151 wl_105 vdd gnd cell_6t
Xbit_r106_c151 bl_151 br_151 wl_106 vdd gnd cell_6t
Xbit_r107_c151 bl_151 br_151 wl_107 vdd gnd cell_6t
Xbit_r108_c151 bl_151 br_151 wl_108 vdd gnd cell_6t
Xbit_r109_c151 bl_151 br_151 wl_109 vdd gnd cell_6t
Xbit_r110_c151 bl_151 br_151 wl_110 vdd gnd cell_6t
Xbit_r111_c151 bl_151 br_151 wl_111 vdd gnd cell_6t
Xbit_r112_c151 bl_151 br_151 wl_112 vdd gnd cell_6t
Xbit_r113_c151 bl_151 br_151 wl_113 vdd gnd cell_6t
Xbit_r114_c151 bl_151 br_151 wl_114 vdd gnd cell_6t
Xbit_r115_c151 bl_151 br_151 wl_115 vdd gnd cell_6t
Xbit_r116_c151 bl_151 br_151 wl_116 vdd gnd cell_6t
Xbit_r117_c151 bl_151 br_151 wl_117 vdd gnd cell_6t
Xbit_r118_c151 bl_151 br_151 wl_118 vdd gnd cell_6t
Xbit_r119_c151 bl_151 br_151 wl_119 vdd gnd cell_6t
Xbit_r120_c151 bl_151 br_151 wl_120 vdd gnd cell_6t
Xbit_r121_c151 bl_151 br_151 wl_121 vdd gnd cell_6t
Xbit_r122_c151 bl_151 br_151 wl_122 vdd gnd cell_6t
Xbit_r123_c151 bl_151 br_151 wl_123 vdd gnd cell_6t
Xbit_r124_c151 bl_151 br_151 wl_124 vdd gnd cell_6t
Xbit_r125_c151 bl_151 br_151 wl_125 vdd gnd cell_6t
Xbit_r126_c151 bl_151 br_151 wl_126 vdd gnd cell_6t
Xbit_r127_c151 bl_151 br_151 wl_127 vdd gnd cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd cell_6t
Xbit_r1_c152 bl_152 br_152 wl_1 vdd gnd cell_6t
Xbit_r2_c152 bl_152 br_152 wl_2 vdd gnd cell_6t
Xbit_r3_c152 bl_152 br_152 wl_3 vdd gnd cell_6t
Xbit_r4_c152 bl_152 br_152 wl_4 vdd gnd cell_6t
Xbit_r5_c152 bl_152 br_152 wl_5 vdd gnd cell_6t
Xbit_r6_c152 bl_152 br_152 wl_6 vdd gnd cell_6t
Xbit_r7_c152 bl_152 br_152 wl_7 vdd gnd cell_6t
Xbit_r8_c152 bl_152 br_152 wl_8 vdd gnd cell_6t
Xbit_r9_c152 bl_152 br_152 wl_9 vdd gnd cell_6t
Xbit_r10_c152 bl_152 br_152 wl_10 vdd gnd cell_6t
Xbit_r11_c152 bl_152 br_152 wl_11 vdd gnd cell_6t
Xbit_r12_c152 bl_152 br_152 wl_12 vdd gnd cell_6t
Xbit_r13_c152 bl_152 br_152 wl_13 vdd gnd cell_6t
Xbit_r14_c152 bl_152 br_152 wl_14 vdd gnd cell_6t
Xbit_r15_c152 bl_152 br_152 wl_15 vdd gnd cell_6t
Xbit_r16_c152 bl_152 br_152 wl_16 vdd gnd cell_6t
Xbit_r17_c152 bl_152 br_152 wl_17 vdd gnd cell_6t
Xbit_r18_c152 bl_152 br_152 wl_18 vdd gnd cell_6t
Xbit_r19_c152 bl_152 br_152 wl_19 vdd gnd cell_6t
Xbit_r20_c152 bl_152 br_152 wl_20 vdd gnd cell_6t
Xbit_r21_c152 bl_152 br_152 wl_21 vdd gnd cell_6t
Xbit_r22_c152 bl_152 br_152 wl_22 vdd gnd cell_6t
Xbit_r23_c152 bl_152 br_152 wl_23 vdd gnd cell_6t
Xbit_r24_c152 bl_152 br_152 wl_24 vdd gnd cell_6t
Xbit_r25_c152 bl_152 br_152 wl_25 vdd gnd cell_6t
Xbit_r26_c152 bl_152 br_152 wl_26 vdd gnd cell_6t
Xbit_r27_c152 bl_152 br_152 wl_27 vdd gnd cell_6t
Xbit_r28_c152 bl_152 br_152 wl_28 vdd gnd cell_6t
Xbit_r29_c152 bl_152 br_152 wl_29 vdd gnd cell_6t
Xbit_r30_c152 bl_152 br_152 wl_30 vdd gnd cell_6t
Xbit_r31_c152 bl_152 br_152 wl_31 vdd gnd cell_6t
Xbit_r32_c152 bl_152 br_152 wl_32 vdd gnd cell_6t
Xbit_r33_c152 bl_152 br_152 wl_33 vdd gnd cell_6t
Xbit_r34_c152 bl_152 br_152 wl_34 vdd gnd cell_6t
Xbit_r35_c152 bl_152 br_152 wl_35 vdd gnd cell_6t
Xbit_r36_c152 bl_152 br_152 wl_36 vdd gnd cell_6t
Xbit_r37_c152 bl_152 br_152 wl_37 vdd gnd cell_6t
Xbit_r38_c152 bl_152 br_152 wl_38 vdd gnd cell_6t
Xbit_r39_c152 bl_152 br_152 wl_39 vdd gnd cell_6t
Xbit_r40_c152 bl_152 br_152 wl_40 vdd gnd cell_6t
Xbit_r41_c152 bl_152 br_152 wl_41 vdd gnd cell_6t
Xbit_r42_c152 bl_152 br_152 wl_42 vdd gnd cell_6t
Xbit_r43_c152 bl_152 br_152 wl_43 vdd gnd cell_6t
Xbit_r44_c152 bl_152 br_152 wl_44 vdd gnd cell_6t
Xbit_r45_c152 bl_152 br_152 wl_45 vdd gnd cell_6t
Xbit_r46_c152 bl_152 br_152 wl_46 vdd gnd cell_6t
Xbit_r47_c152 bl_152 br_152 wl_47 vdd gnd cell_6t
Xbit_r48_c152 bl_152 br_152 wl_48 vdd gnd cell_6t
Xbit_r49_c152 bl_152 br_152 wl_49 vdd gnd cell_6t
Xbit_r50_c152 bl_152 br_152 wl_50 vdd gnd cell_6t
Xbit_r51_c152 bl_152 br_152 wl_51 vdd gnd cell_6t
Xbit_r52_c152 bl_152 br_152 wl_52 vdd gnd cell_6t
Xbit_r53_c152 bl_152 br_152 wl_53 vdd gnd cell_6t
Xbit_r54_c152 bl_152 br_152 wl_54 vdd gnd cell_6t
Xbit_r55_c152 bl_152 br_152 wl_55 vdd gnd cell_6t
Xbit_r56_c152 bl_152 br_152 wl_56 vdd gnd cell_6t
Xbit_r57_c152 bl_152 br_152 wl_57 vdd gnd cell_6t
Xbit_r58_c152 bl_152 br_152 wl_58 vdd gnd cell_6t
Xbit_r59_c152 bl_152 br_152 wl_59 vdd gnd cell_6t
Xbit_r60_c152 bl_152 br_152 wl_60 vdd gnd cell_6t
Xbit_r61_c152 bl_152 br_152 wl_61 vdd gnd cell_6t
Xbit_r62_c152 bl_152 br_152 wl_62 vdd gnd cell_6t
Xbit_r63_c152 bl_152 br_152 wl_63 vdd gnd cell_6t
Xbit_r64_c152 bl_152 br_152 wl_64 vdd gnd cell_6t
Xbit_r65_c152 bl_152 br_152 wl_65 vdd gnd cell_6t
Xbit_r66_c152 bl_152 br_152 wl_66 vdd gnd cell_6t
Xbit_r67_c152 bl_152 br_152 wl_67 vdd gnd cell_6t
Xbit_r68_c152 bl_152 br_152 wl_68 vdd gnd cell_6t
Xbit_r69_c152 bl_152 br_152 wl_69 vdd gnd cell_6t
Xbit_r70_c152 bl_152 br_152 wl_70 vdd gnd cell_6t
Xbit_r71_c152 bl_152 br_152 wl_71 vdd gnd cell_6t
Xbit_r72_c152 bl_152 br_152 wl_72 vdd gnd cell_6t
Xbit_r73_c152 bl_152 br_152 wl_73 vdd gnd cell_6t
Xbit_r74_c152 bl_152 br_152 wl_74 vdd gnd cell_6t
Xbit_r75_c152 bl_152 br_152 wl_75 vdd gnd cell_6t
Xbit_r76_c152 bl_152 br_152 wl_76 vdd gnd cell_6t
Xbit_r77_c152 bl_152 br_152 wl_77 vdd gnd cell_6t
Xbit_r78_c152 bl_152 br_152 wl_78 vdd gnd cell_6t
Xbit_r79_c152 bl_152 br_152 wl_79 vdd gnd cell_6t
Xbit_r80_c152 bl_152 br_152 wl_80 vdd gnd cell_6t
Xbit_r81_c152 bl_152 br_152 wl_81 vdd gnd cell_6t
Xbit_r82_c152 bl_152 br_152 wl_82 vdd gnd cell_6t
Xbit_r83_c152 bl_152 br_152 wl_83 vdd gnd cell_6t
Xbit_r84_c152 bl_152 br_152 wl_84 vdd gnd cell_6t
Xbit_r85_c152 bl_152 br_152 wl_85 vdd gnd cell_6t
Xbit_r86_c152 bl_152 br_152 wl_86 vdd gnd cell_6t
Xbit_r87_c152 bl_152 br_152 wl_87 vdd gnd cell_6t
Xbit_r88_c152 bl_152 br_152 wl_88 vdd gnd cell_6t
Xbit_r89_c152 bl_152 br_152 wl_89 vdd gnd cell_6t
Xbit_r90_c152 bl_152 br_152 wl_90 vdd gnd cell_6t
Xbit_r91_c152 bl_152 br_152 wl_91 vdd gnd cell_6t
Xbit_r92_c152 bl_152 br_152 wl_92 vdd gnd cell_6t
Xbit_r93_c152 bl_152 br_152 wl_93 vdd gnd cell_6t
Xbit_r94_c152 bl_152 br_152 wl_94 vdd gnd cell_6t
Xbit_r95_c152 bl_152 br_152 wl_95 vdd gnd cell_6t
Xbit_r96_c152 bl_152 br_152 wl_96 vdd gnd cell_6t
Xbit_r97_c152 bl_152 br_152 wl_97 vdd gnd cell_6t
Xbit_r98_c152 bl_152 br_152 wl_98 vdd gnd cell_6t
Xbit_r99_c152 bl_152 br_152 wl_99 vdd gnd cell_6t
Xbit_r100_c152 bl_152 br_152 wl_100 vdd gnd cell_6t
Xbit_r101_c152 bl_152 br_152 wl_101 vdd gnd cell_6t
Xbit_r102_c152 bl_152 br_152 wl_102 vdd gnd cell_6t
Xbit_r103_c152 bl_152 br_152 wl_103 vdd gnd cell_6t
Xbit_r104_c152 bl_152 br_152 wl_104 vdd gnd cell_6t
Xbit_r105_c152 bl_152 br_152 wl_105 vdd gnd cell_6t
Xbit_r106_c152 bl_152 br_152 wl_106 vdd gnd cell_6t
Xbit_r107_c152 bl_152 br_152 wl_107 vdd gnd cell_6t
Xbit_r108_c152 bl_152 br_152 wl_108 vdd gnd cell_6t
Xbit_r109_c152 bl_152 br_152 wl_109 vdd gnd cell_6t
Xbit_r110_c152 bl_152 br_152 wl_110 vdd gnd cell_6t
Xbit_r111_c152 bl_152 br_152 wl_111 vdd gnd cell_6t
Xbit_r112_c152 bl_152 br_152 wl_112 vdd gnd cell_6t
Xbit_r113_c152 bl_152 br_152 wl_113 vdd gnd cell_6t
Xbit_r114_c152 bl_152 br_152 wl_114 vdd gnd cell_6t
Xbit_r115_c152 bl_152 br_152 wl_115 vdd gnd cell_6t
Xbit_r116_c152 bl_152 br_152 wl_116 vdd gnd cell_6t
Xbit_r117_c152 bl_152 br_152 wl_117 vdd gnd cell_6t
Xbit_r118_c152 bl_152 br_152 wl_118 vdd gnd cell_6t
Xbit_r119_c152 bl_152 br_152 wl_119 vdd gnd cell_6t
Xbit_r120_c152 bl_152 br_152 wl_120 vdd gnd cell_6t
Xbit_r121_c152 bl_152 br_152 wl_121 vdd gnd cell_6t
Xbit_r122_c152 bl_152 br_152 wl_122 vdd gnd cell_6t
Xbit_r123_c152 bl_152 br_152 wl_123 vdd gnd cell_6t
Xbit_r124_c152 bl_152 br_152 wl_124 vdd gnd cell_6t
Xbit_r125_c152 bl_152 br_152 wl_125 vdd gnd cell_6t
Xbit_r126_c152 bl_152 br_152 wl_126 vdd gnd cell_6t
Xbit_r127_c152 bl_152 br_152 wl_127 vdd gnd cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd cell_6t
Xbit_r1_c153 bl_153 br_153 wl_1 vdd gnd cell_6t
Xbit_r2_c153 bl_153 br_153 wl_2 vdd gnd cell_6t
Xbit_r3_c153 bl_153 br_153 wl_3 vdd gnd cell_6t
Xbit_r4_c153 bl_153 br_153 wl_4 vdd gnd cell_6t
Xbit_r5_c153 bl_153 br_153 wl_5 vdd gnd cell_6t
Xbit_r6_c153 bl_153 br_153 wl_6 vdd gnd cell_6t
Xbit_r7_c153 bl_153 br_153 wl_7 vdd gnd cell_6t
Xbit_r8_c153 bl_153 br_153 wl_8 vdd gnd cell_6t
Xbit_r9_c153 bl_153 br_153 wl_9 vdd gnd cell_6t
Xbit_r10_c153 bl_153 br_153 wl_10 vdd gnd cell_6t
Xbit_r11_c153 bl_153 br_153 wl_11 vdd gnd cell_6t
Xbit_r12_c153 bl_153 br_153 wl_12 vdd gnd cell_6t
Xbit_r13_c153 bl_153 br_153 wl_13 vdd gnd cell_6t
Xbit_r14_c153 bl_153 br_153 wl_14 vdd gnd cell_6t
Xbit_r15_c153 bl_153 br_153 wl_15 vdd gnd cell_6t
Xbit_r16_c153 bl_153 br_153 wl_16 vdd gnd cell_6t
Xbit_r17_c153 bl_153 br_153 wl_17 vdd gnd cell_6t
Xbit_r18_c153 bl_153 br_153 wl_18 vdd gnd cell_6t
Xbit_r19_c153 bl_153 br_153 wl_19 vdd gnd cell_6t
Xbit_r20_c153 bl_153 br_153 wl_20 vdd gnd cell_6t
Xbit_r21_c153 bl_153 br_153 wl_21 vdd gnd cell_6t
Xbit_r22_c153 bl_153 br_153 wl_22 vdd gnd cell_6t
Xbit_r23_c153 bl_153 br_153 wl_23 vdd gnd cell_6t
Xbit_r24_c153 bl_153 br_153 wl_24 vdd gnd cell_6t
Xbit_r25_c153 bl_153 br_153 wl_25 vdd gnd cell_6t
Xbit_r26_c153 bl_153 br_153 wl_26 vdd gnd cell_6t
Xbit_r27_c153 bl_153 br_153 wl_27 vdd gnd cell_6t
Xbit_r28_c153 bl_153 br_153 wl_28 vdd gnd cell_6t
Xbit_r29_c153 bl_153 br_153 wl_29 vdd gnd cell_6t
Xbit_r30_c153 bl_153 br_153 wl_30 vdd gnd cell_6t
Xbit_r31_c153 bl_153 br_153 wl_31 vdd gnd cell_6t
Xbit_r32_c153 bl_153 br_153 wl_32 vdd gnd cell_6t
Xbit_r33_c153 bl_153 br_153 wl_33 vdd gnd cell_6t
Xbit_r34_c153 bl_153 br_153 wl_34 vdd gnd cell_6t
Xbit_r35_c153 bl_153 br_153 wl_35 vdd gnd cell_6t
Xbit_r36_c153 bl_153 br_153 wl_36 vdd gnd cell_6t
Xbit_r37_c153 bl_153 br_153 wl_37 vdd gnd cell_6t
Xbit_r38_c153 bl_153 br_153 wl_38 vdd gnd cell_6t
Xbit_r39_c153 bl_153 br_153 wl_39 vdd gnd cell_6t
Xbit_r40_c153 bl_153 br_153 wl_40 vdd gnd cell_6t
Xbit_r41_c153 bl_153 br_153 wl_41 vdd gnd cell_6t
Xbit_r42_c153 bl_153 br_153 wl_42 vdd gnd cell_6t
Xbit_r43_c153 bl_153 br_153 wl_43 vdd gnd cell_6t
Xbit_r44_c153 bl_153 br_153 wl_44 vdd gnd cell_6t
Xbit_r45_c153 bl_153 br_153 wl_45 vdd gnd cell_6t
Xbit_r46_c153 bl_153 br_153 wl_46 vdd gnd cell_6t
Xbit_r47_c153 bl_153 br_153 wl_47 vdd gnd cell_6t
Xbit_r48_c153 bl_153 br_153 wl_48 vdd gnd cell_6t
Xbit_r49_c153 bl_153 br_153 wl_49 vdd gnd cell_6t
Xbit_r50_c153 bl_153 br_153 wl_50 vdd gnd cell_6t
Xbit_r51_c153 bl_153 br_153 wl_51 vdd gnd cell_6t
Xbit_r52_c153 bl_153 br_153 wl_52 vdd gnd cell_6t
Xbit_r53_c153 bl_153 br_153 wl_53 vdd gnd cell_6t
Xbit_r54_c153 bl_153 br_153 wl_54 vdd gnd cell_6t
Xbit_r55_c153 bl_153 br_153 wl_55 vdd gnd cell_6t
Xbit_r56_c153 bl_153 br_153 wl_56 vdd gnd cell_6t
Xbit_r57_c153 bl_153 br_153 wl_57 vdd gnd cell_6t
Xbit_r58_c153 bl_153 br_153 wl_58 vdd gnd cell_6t
Xbit_r59_c153 bl_153 br_153 wl_59 vdd gnd cell_6t
Xbit_r60_c153 bl_153 br_153 wl_60 vdd gnd cell_6t
Xbit_r61_c153 bl_153 br_153 wl_61 vdd gnd cell_6t
Xbit_r62_c153 bl_153 br_153 wl_62 vdd gnd cell_6t
Xbit_r63_c153 bl_153 br_153 wl_63 vdd gnd cell_6t
Xbit_r64_c153 bl_153 br_153 wl_64 vdd gnd cell_6t
Xbit_r65_c153 bl_153 br_153 wl_65 vdd gnd cell_6t
Xbit_r66_c153 bl_153 br_153 wl_66 vdd gnd cell_6t
Xbit_r67_c153 bl_153 br_153 wl_67 vdd gnd cell_6t
Xbit_r68_c153 bl_153 br_153 wl_68 vdd gnd cell_6t
Xbit_r69_c153 bl_153 br_153 wl_69 vdd gnd cell_6t
Xbit_r70_c153 bl_153 br_153 wl_70 vdd gnd cell_6t
Xbit_r71_c153 bl_153 br_153 wl_71 vdd gnd cell_6t
Xbit_r72_c153 bl_153 br_153 wl_72 vdd gnd cell_6t
Xbit_r73_c153 bl_153 br_153 wl_73 vdd gnd cell_6t
Xbit_r74_c153 bl_153 br_153 wl_74 vdd gnd cell_6t
Xbit_r75_c153 bl_153 br_153 wl_75 vdd gnd cell_6t
Xbit_r76_c153 bl_153 br_153 wl_76 vdd gnd cell_6t
Xbit_r77_c153 bl_153 br_153 wl_77 vdd gnd cell_6t
Xbit_r78_c153 bl_153 br_153 wl_78 vdd gnd cell_6t
Xbit_r79_c153 bl_153 br_153 wl_79 vdd gnd cell_6t
Xbit_r80_c153 bl_153 br_153 wl_80 vdd gnd cell_6t
Xbit_r81_c153 bl_153 br_153 wl_81 vdd gnd cell_6t
Xbit_r82_c153 bl_153 br_153 wl_82 vdd gnd cell_6t
Xbit_r83_c153 bl_153 br_153 wl_83 vdd gnd cell_6t
Xbit_r84_c153 bl_153 br_153 wl_84 vdd gnd cell_6t
Xbit_r85_c153 bl_153 br_153 wl_85 vdd gnd cell_6t
Xbit_r86_c153 bl_153 br_153 wl_86 vdd gnd cell_6t
Xbit_r87_c153 bl_153 br_153 wl_87 vdd gnd cell_6t
Xbit_r88_c153 bl_153 br_153 wl_88 vdd gnd cell_6t
Xbit_r89_c153 bl_153 br_153 wl_89 vdd gnd cell_6t
Xbit_r90_c153 bl_153 br_153 wl_90 vdd gnd cell_6t
Xbit_r91_c153 bl_153 br_153 wl_91 vdd gnd cell_6t
Xbit_r92_c153 bl_153 br_153 wl_92 vdd gnd cell_6t
Xbit_r93_c153 bl_153 br_153 wl_93 vdd gnd cell_6t
Xbit_r94_c153 bl_153 br_153 wl_94 vdd gnd cell_6t
Xbit_r95_c153 bl_153 br_153 wl_95 vdd gnd cell_6t
Xbit_r96_c153 bl_153 br_153 wl_96 vdd gnd cell_6t
Xbit_r97_c153 bl_153 br_153 wl_97 vdd gnd cell_6t
Xbit_r98_c153 bl_153 br_153 wl_98 vdd gnd cell_6t
Xbit_r99_c153 bl_153 br_153 wl_99 vdd gnd cell_6t
Xbit_r100_c153 bl_153 br_153 wl_100 vdd gnd cell_6t
Xbit_r101_c153 bl_153 br_153 wl_101 vdd gnd cell_6t
Xbit_r102_c153 bl_153 br_153 wl_102 vdd gnd cell_6t
Xbit_r103_c153 bl_153 br_153 wl_103 vdd gnd cell_6t
Xbit_r104_c153 bl_153 br_153 wl_104 vdd gnd cell_6t
Xbit_r105_c153 bl_153 br_153 wl_105 vdd gnd cell_6t
Xbit_r106_c153 bl_153 br_153 wl_106 vdd gnd cell_6t
Xbit_r107_c153 bl_153 br_153 wl_107 vdd gnd cell_6t
Xbit_r108_c153 bl_153 br_153 wl_108 vdd gnd cell_6t
Xbit_r109_c153 bl_153 br_153 wl_109 vdd gnd cell_6t
Xbit_r110_c153 bl_153 br_153 wl_110 vdd gnd cell_6t
Xbit_r111_c153 bl_153 br_153 wl_111 vdd gnd cell_6t
Xbit_r112_c153 bl_153 br_153 wl_112 vdd gnd cell_6t
Xbit_r113_c153 bl_153 br_153 wl_113 vdd gnd cell_6t
Xbit_r114_c153 bl_153 br_153 wl_114 vdd gnd cell_6t
Xbit_r115_c153 bl_153 br_153 wl_115 vdd gnd cell_6t
Xbit_r116_c153 bl_153 br_153 wl_116 vdd gnd cell_6t
Xbit_r117_c153 bl_153 br_153 wl_117 vdd gnd cell_6t
Xbit_r118_c153 bl_153 br_153 wl_118 vdd gnd cell_6t
Xbit_r119_c153 bl_153 br_153 wl_119 vdd gnd cell_6t
Xbit_r120_c153 bl_153 br_153 wl_120 vdd gnd cell_6t
Xbit_r121_c153 bl_153 br_153 wl_121 vdd gnd cell_6t
Xbit_r122_c153 bl_153 br_153 wl_122 vdd gnd cell_6t
Xbit_r123_c153 bl_153 br_153 wl_123 vdd gnd cell_6t
Xbit_r124_c153 bl_153 br_153 wl_124 vdd gnd cell_6t
Xbit_r125_c153 bl_153 br_153 wl_125 vdd gnd cell_6t
Xbit_r126_c153 bl_153 br_153 wl_126 vdd gnd cell_6t
Xbit_r127_c153 bl_153 br_153 wl_127 vdd gnd cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd cell_6t
Xbit_r1_c154 bl_154 br_154 wl_1 vdd gnd cell_6t
Xbit_r2_c154 bl_154 br_154 wl_2 vdd gnd cell_6t
Xbit_r3_c154 bl_154 br_154 wl_3 vdd gnd cell_6t
Xbit_r4_c154 bl_154 br_154 wl_4 vdd gnd cell_6t
Xbit_r5_c154 bl_154 br_154 wl_5 vdd gnd cell_6t
Xbit_r6_c154 bl_154 br_154 wl_6 vdd gnd cell_6t
Xbit_r7_c154 bl_154 br_154 wl_7 vdd gnd cell_6t
Xbit_r8_c154 bl_154 br_154 wl_8 vdd gnd cell_6t
Xbit_r9_c154 bl_154 br_154 wl_9 vdd gnd cell_6t
Xbit_r10_c154 bl_154 br_154 wl_10 vdd gnd cell_6t
Xbit_r11_c154 bl_154 br_154 wl_11 vdd gnd cell_6t
Xbit_r12_c154 bl_154 br_154 wl_12 vdd gnd cell_6t
Xbit_r13_c154 bl_154 br_154 wl_13 vdd gnd cell_6t
Xbit_r14_c154 bl_154 br_154 wl_14 vdd gnd cell_6t
Xbit_r15_c154 bl_154 br_154 wl_15 vdd gnd cell_6t
Xbit_r16_c154 bl_154 br_154 wl_16 vdd gnd cell_6t
Xbit_r17_c154 bl_154 br_154 wl_17 vdd gnd cell_6t
Xbit_r18_c154 bl_154 br_154 wl_18 vdd gnd cell_6t
Xbit_r19_c154 bl_154 br_154 wl_19 vdd gnd cell_6t
Xbit_r20_c154 bl_154 br_154 wl_20 vdd gnd cell_6t
Xbit_r21_c154 bl_154 br_154 wl_21 vdd gnd cell_6t
Xbit_r22_c154 bl_154 br_154 wl_22 vdd gnd cell_6t
Xbit_r23_c154 bl_154 br_154 wl_23 vdd gnd cell_6t
Xbit_r24_c154 bl_154 br_154 wl_24 vdd gnd cell_6t
Xbit_r25_c154 bl_154 br_154 wl_25 vdd gnd cell_6t
Xbit_r26_c154 bl_154 br_154 wl_26 vdd gnd cell_6t
Xbit_r27_c154 bl_154 br_154 wl_27 vdd gnd cell_6t
Xbit_r28_c154 bl_154 br_154 wl_28 vdd gnd cell_6t
Xbit_r29_c154 bl_154 br_154 wl_29 vdd gnd cell_6t
Xbit_r30_c154 bl_154 br_154 wl_30 vdd gnd cell_6t
Xbit_r31_c154 bl_154 br_154 wl_31 vdd gnd cell_6t
Xbit_r32_c154 bl_154 br_154 wl_32 vdd gnd cell_6t
Xbit_r33_c154 bl_154 br_154 wl_33 vdd gnd cell_6t
Xbit_r34_c154 bl_154 br_154 wl_34 vdd gnd cell_6t
Xbit_r35_c154 bl_154 br_154 wl_35 vdd gnd cell_6t
Xbit_r36_c154 bl_154 br_154 wl_36 vdd gnd cell_6t
Xbit_r37_c154 bl_154 br_154 wl_37 vdd gnd cell_6t
Xbit_r38_c154 bl_154 br_154 wl_38 vdd gnd cell_6t
Xbit_r39_c154 bl_154 br_154 wl_39 vdd gnd cell_6t
Xbit_r40_c154 bl_154 br_154 wl_40 vdd gnd cell_6t
Xbit_r41_c154 bl_154 br_154 wl_41 vdd gnd cell_6t
Xbit_r42_c154 bl_154 br_154 wl_42 vdd gnd cell_6t
Xbit_r43_c154 bl_154 br_154 wl_43 vdd gnd cell_6t
Xbit_r44_c154 bl_154 br_154 wl_44 vdd gnd cell_6t
Xbit_r45_c154 bl_154 br_154 wl_45 vdd gnd cell_6t
Xbit_r46_c154 bl_154 br_154 wl_46 vdd gnd cell_6t
Xbit_r47_c154 bl_154 br_154 wl_47 vdd gnd cell_6t
Xbit_r48_c154 bl_154 br_154 wl_48 vdd gnd cell_6t
Xbit_r49_c154 bl_154 br_154 wl_49 vdd gnd cell_6t
Xbit_r50_c154 bl_154 br_154 wl_50 vdd gnd cell_6t
Xbit_r51_c154 bl_154 br_154 wl_51 vdd gnd cell_6t
Xbit_r52_c154 bl_154 br_154 wl_52 vdd gnd cell_6t
Xbit_r53_c154 bl_154 br_154 wl_53 vdd gnd cell_6t
Xbit_r54_c154 bl_154 br_154 wl_54 vdd gnd cell_6t
Xbit_r55_c154 bl_154 br_154 wl_55 vdd gnd cell_6t
Xbit_r56_c154 bl_154 br_154 wl_56 vdd gnd cell_6t
Xbit_r57_c154 bl_154 br_154 wl_57 vdd gnd cell_6t
Xbit_r58_c154 bl_154 br_154 wl_58 vdd gnd cell_6t
Xbit_r59_c154 bl_154 br_154 wl_59 vdd gnd cell_6t
Xbit_r60_c154 bl_154 br_154 wl_60 vdd gnd cell_6t
Xbit_r61_c154 bl_154 br_154 wl_61 vdd gnd cell_6t
Xbit_r62_c154 bl_154 br_154 wl_62 vdd gnd cell_6t
Xbit_r63_c154 bl_154 br_154 wl_63 vdd gnd cell_6t
Xbit_r64_c154 bl_154 br_154 wl_64 vdd gnd cell_6t
Xbit_r65_c154 bl_154 br_154 wl_65 vdd gnd cell_6t
Xbit_r66_c154 bl_154 br_154 wl_66 vdd gnd cell_6t
Xbit_r67_c154 bl_154 br_154 wl_67 vdd gnd cell_6t
Xbit_r68_c154 bl_154 br_154 wl_68 vdd gnd cell_6t
Xbit_r69_c154 bl_154 br_154 wl_69 vdd gnd cell_6t
Xbit_r70_c154 bl_154 br_154 wl_70 vdd gnd cell_6t
Xbit_r71_c154 bl_154 br_154 wl_71 vdd gnd cell_6t
Xbit_r72_c154 bl_154 br_154 wl_72 vdd gnd cell_6t
Xbit_r73_c154 bl_154 br_154 wl_73 vdd gnd cell_6t
Xbit_r74_c154 bl_154 br_154 wl_74 vdd gnd cell_6t
Xbit_r75_c154 bl_154 br_154 wl_75 vdd gnd cell_6t
Xbit_r76_c154 bl_154 br_154 wl_76 vdd gnd cell_6t
Xbit_r77_c154 bl_154 br_154 wl_77 vdd gnd cell_6t
Xbit_r78_c154 bl_154 br_154 wl_78 vdd gnd cell_6t
Xbit_r79_c154 bl_154 br_154 wl_79 vdd gnd cell_6t
Xbit_r80_c154 bl_154 br_154 wl_80 vdd gnd cell_6t
Xbit_r81_c154 bl_154 br_154 wl_81 vdd gnd cell_6t
Xbit_r82_c154 bl_154 br_154 wl_82 vdd gnd cell_6t
Xbit_r83_c154 bl_154 br_154 wl_83 vdd gnd cell_6t
Xbit_r84_c154 bl_154 br_154 wl_84 vdd gnd cell_6t
Xbit_r85_c154 bl_154 br_154 wl_85 vdd gnd cell_6t
Xbit_r86_c154 bl_154 br_154 wl_86 vdd gnd cell_6t
Xbit_r87_c154 bl_154 br_154 wl_87 vdd gnd cell_6t
Xbit_r88_c154 bl_154 br_154 wl_88 vdd gnd cell_6t
Xbit_r89_c154 bl_154 br_154 wl_89 vdd gnd cell_6t
Xbit_r90_c154 bl_154 br_154 wl_90 vdd gnd cell_6t
Xbit_r91_c154 bl_154 br_154 wl_91 vdd gnd cell_6t
Xbit_r92_c154 bl_154 br_154 wl_92 vdd gnd cell_6t
Xbit_r93_c154 bl_154 br_154 wl_93 vdd gnd cell_6t
Xbit_r94_c154 bl_154 br_154 wl_94 vdd gnd cell_6t
Xbit_r95_c154 bl_154 br_154 wl_95 vdd gnd cell_6t
Xbit_r96_c154 bl_154 br_154 wl_96 vdd gnd cell_6t
Xbit_r97_c154 bl_154 br_154 wl_97 vdd gnd cell_6t
Xbit_r98_c154 bl_154 br_154 wl_98 vdd gnd cell_6t
Xbit_r99_c154 bl_154 br_154 wl_99 vdd gnd cell_6t
Xbit_r100_c154 bl_154 br_154 wl_100 vdd gnd cell_6t
Xbit_r101_c154 bl_154 br_154 wl_101 vdd gnd cell_6t
Xbit_r102_c154 bl_154 br_154 wl_102 vdd gnd cell_6t
Xbit_r103_c154 bl_154 br_154 wl_103 vdd gnd cell_6t
Xbit_r104_c154 bl_154 br_154 wl_104 vdd gnd cell_6t
Xbit_r105_c154 bl_154 br_154 wl_105 vdd gnd cell_6t
Xbit_r106_c154 bl_154 br_154 wl_106 vdd gnd cell_6t
Xbit_r107_c154 bl_154 br_154 wl_107 vdd gnd cell_6t
Xbit_r108_c154 bl_154 br_154 wl_108 vdd gnd cell_6t
Xbit_r109_c154 bl_154 br_154 wl_109 vdd gnd cell_6t
Xbit_r110_c154 bl_154 br_154 wl_110 vdd gnd cell_6t
Xbit_r111_c154 bl_154 br_154 wl_111 vdd gnd cell_6t
Xbit_r112_c154 bl_154 br_154 wl_112 vdd gnd cell_6t
Xbit_r113_c154 bl_154 br_154 wl_113 vdd gnd cell_6t
Xbit_r114_c154 bl_154 br_154 wl_114 vdd gnd cell_6t
Xbit_r115_c154 bl_154 br_154 wl_115 vdd gnd cell_6t
Xbit_r116_c154 bl_154 br_154 wl_116 vdd gnd cell_6t
Xbit_r117_c154 bl_154 br_154 wl_117 vdd gnd cell_6t
Xbit_r118_c154 bl_154 br_154 wl_118 vdd gnd cell_6t
Xbit_r119_c154 bl_154 br_154 wl_119 vdd gnd cell_6t
Xbit_r120_c154 bl_154 br_154 wl_120 vdd gnd cell_6t
Xbit_r121_c154 bl_154 br_154 wl_121 vdd gnd cell_6t
Xbit_r122_c154 bl_154 br_154 wl_122 vdd gnd cell_6t
Xbit_r123_c154 bl_154 br_154 wl_123 vdd gnd cell_6t
Xbit_r124_c154 bl_154 br_154 wl_124 vdd gnd cell_6t
Xbit_r125_c154 bl_154 br_154 wl_125 vdd gnd cell_6t
Xbit_r126_c154 bl_154 br_154 wl_126 vdd gnd cell_6t
Xbit_r127_c154 bl_154 br_154 wl_127 vdd gnd cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd cell_6t
Xbit_r1_c155 bl_155 br_155 wl_1 vdd gnd cell_6t
Xbit_r2_c155 bl_155 br_155 wl_2 vdd gnd cell_6t
Xbit_r3_c155 bl_155 br_155 wl_3 vdd gnd cell_6t
Xbit_r4_c155 bl_155 br_155 wl_4 vdd gnd cell_6t
Xbit_r5_c155 bl_155 br_155 wl_5 vdd gnd cell_6t
Xbit_r6_c155 bl_155 br_155 wl_6 vdd gnd cell_6t
Xbit_r7_c155 bl_155 br_155 wl_7 vdd gnd cell_6t
Xbit_r8_c155 bl_155 br_155 wl_8 vdd gnd cell_6t
Xbit_r9_c155 bl_155 br_155 wl_9 vdd gnd cell_6t
Xbit_r10_c155 bl_155 br_155 wl_10 vdd gnd cell_6t
Xbit_r11_c155 bl_155 br_155 wl_11 vdd gnd cell_6t
Xbit_r12_c155 bl_155 br_155 wl_12 vdd gnd cell_6t
Xbit_r13_c155 bl_155 br_155 wl_13 vdd gnd cell_6t
Xbit_r14_c155 bl_155 br_155 wl_14 vdd gnd cell_6t
Xbit_r15_c155 bl_155 br_155 wl_15 vdd gnd cell_6t
Xbit_r16_c155 bl_155 br_155 wl_16 vdd gnd cell_6t
Xbit_r17_c155 bl_155 br_155 wl_17 vdd gnd cell_6t
Xbit_r18_c155 bl_155 br_155 wl_18 vdd gnd cell_6t
Xbit_r19_c155 bl_155 br_155 wl_19 vdd gnd cell_6t
Xbit_r20_c155 bl_155 br_155 wl_20 vdd gnd cell_6t
Xbit_r21_c155 bl_155 br_155 wl_21 vdd gnd cell_6t
Xbit_r22_c155 bl_155 br_155 wl_22 vdd gnd cell_6t
Xbit_r23_c155 bl_155 br_155 wl_23 vdd gnd cell_6t
Xbit_r24_c155 bl_155 br_155 wl_24 vdd gnd cell_6t
Xbit_r25_c155 bl_155 br_155 wl_25 vdd gnd cell_6t
Xbit_r26_c155 bl_155 br_155 wl_26 vdd gnd cell_6t
Xbit_r27_c155 bl_155 br_155 wl_27 vdd gnd cell_6t
Xbit_r28_c155 bl_155 br_155 wl_28 vdd gnd cell_6t
Xbit_r29_c155 bl_155 br_155 wl_29 vdd gnd cell_6t
Xbit_r30_c155 bl_155 br_155 wl_30 vdd gnd cell_6t
Xbit_r31_c155 bl_155 br_155 wl_31 vdd gnd cell_6t
Xbit_r32_c155 bl_155 br_155 wl_32 vdd gnd cell_6t
Xbit_r33_c155 bl_155 br_155 wl_33 vdd gnd cell_6t
Xbit_r34_c155 bl_155 br_155 wl_34 vdd gnd cell_6t
Xbit_r35_c155 bl_155 br_155 wl_35 vdd gnd cell_6t
Xbit_r36_c155 bl_155 br_155 wl_36 vdd gnd cell_6t
Xbit_r37_c155 bl_155 br_155 wl_37 vdd gnd cell_6t
Xbit_r38_c155 bl_155 br_155 wl_38 vdd gnd cell_6t
Xbit_r39_c155 bl_155 br_155 wl_39 vdd gnd cell_6t
Xbit_r40_c155 bl_155 br_155 wl_40 vdd gnd cell_6t
Xbit_r41_c155 bl_155 br_155 wl_41 vdd gnd cell_6t
Xbit_r42_c155 bl_155 br_155 wl_42 vdd gnd cell_6t
Xbit_r43_c155 bl_155 br_155 wl_43 vdd gnd cell_6t
Xbit_r44_c155 bl_155 br_155 wl_44 vdd gnd cell_6t
Xbit_r45_c155 bl_155 br_155 wl_45 vdd gnd cell_6t
Xbit_r46_c155 bl_155 br_155 wl_46 vdd gnd cell_6t
Xbit_r47_c155 bl_155 br_155 wl_47 vdd gnd cell_6t
Xbit_r48_c155 bl_155 br_155 wl_48 vdd gnd cell_6t
Xbit_r49_c155 bl_155 br_155 wl_49 vdd gnd cell_6t
Xbit_r50_c155 bl_155 br_155 wl_50 vdd gnd cell_6t
Xbit_r51_c155 bl_155 br_155 wl_51 vdd gnd cell_6t
Xbit_r52_c155 bl_155 br_155 wl_52 vdd gnd cell_6t
Xbit_r53_c155 bl_155 br_155 wl_53 vdd gnd cell_6t
Xbit_r54_c155 bl_155 br_155 wl_54 vdd gnd cell_6t
Xbit_r55_c155 bl_155 br_155 wl_55 vdd gnd cell_6t
Xbit_r56_c155 bl_155 br_155 wl_56 vdd gnd cell_6t
Xbit_r57_c155 bl_155 br_155 wl_57 vdd gnd cell_6t
Xbit_r58_c155 bl_155 br_155 wl_58 vdd gnd cell_6t
Xbit_r59_c155 bl_155 br_155 wl_59 vdd gnd cell_6t
Xbit_r60_c155 bl_155 br_155 wl_60 vdd gnd cell_6t
Xbit_r61_c155 bl_155 br_155 wl_61 vdd gnd cell_6t
Xbit_r62_c155 bl_155 br_155 wl_62 vdd gnd cell_6t
Xbit_r63_c155 bl_155 br_155 wl_63 vdd gnd cell_6t
Xbit_r64_c155 bl_155 br_155 wl_64 vdd gnd cell_6t
Xbit_r65_c155 bl_155 br_155 wl_65 vdd gnd cell_6t
Xbit_r66_c155 bl_155 br_155 wl_66 vdd gnd cell_6t
Xbit_r67_c155 bl_155 br_155 wl_67 vdd gnd cell_6t
Xbit_r68_c155 bl_155 br_155 wl_68 vdd gnd cell_6t
Xbit_r69_c155 bl_155 br_155 wl_69 vdd gnd cell_6t
Xbit_r70_c155 bl_155 br_155 wl_70 vdd gnd cell_6t
Xbit_r71_c155 bl_155 br_155 wl_71 vdd gnd cell_6t
Xbit_r72_c155 bl_155 br_155 wl_72 vdd gnd cell_6t
Xbit_r73_c155 bl_155 br_155 wl_73 vdd gnd cell_6t
Xbit_r74_c155 bl_155 br_155 wl_74 vdd gnd cell_6t
Xbit_r75_c155 bl_155 br_155 wl_75 vdd gnd cell_6t
Xbit_r76_c155 bl_155 br_155 wl_76 vdd gnd cell_6t
Xbit_r77_c155 bl_155 br_155 wl_77 vdd gnd cell_6t
Xbit_r78_c155 bl_155 br_155 wl_78 vdd gnd cell_6t
Xbit_r79_c155 bl_155 br_155 wl_79 vdd gnd cell_6t
Xbit_r80_c155 bl_155 br_155 wl_80 vdd gnd cell_6t
Xbit_r81_c155 bl_155 br_155 wl_81 vdd gnd cell_6t
Xbit_r82_c155 bl_155 br_155 wl_82 vdd gnd cell_6t
Xbit_r83_c155 bl_155 br_155 wl_83 vdd gnd cell_6t
Xbit_r84_c155 bl_155 br_155 wl_84 vdd gnd cell_6t
Xbit_r85_c155 bl_155 br_155 wl_85 vdd gnd cell_6t
Xbit_r86_c155 bl_155 br_155 wl_86 vdd gnd cell_6t
Xbit_r87_c155 bl_155 br_155 wl_87 vdd gnd cell_6t
Xbit_r88_c155 bl_155 br_155 wl_88 vdd gnd cell_6t
Xbit_r89_c155 bl_155 br_155 wl_89 vdd gnd cell_6t
Xbit_r90_c155 bl_155 br_155 wl_90 vdd gnd cell_6t
Xbit_r91_c155 bl_155 br_155 wl_91 vdd gnd cell_6t
Xbit_r92_c155 bl_155 br_155 wl_92 vdd gnd cell_6t
Xbit_r93_c155 bl_155 br_155 wl_93 vdd gnd cell_6t
Xbit_r94_c155 bl_155 br_155 wl_94 vdd gnd cell_6t
Xbit_r95_c155 bl_155 br_155 wl_95 vdd gnd cell_6t
Xbit_r96_c155 bl_155 br_155 wl_96 vdd gnd cell_6t
Xbit_r97_c155 bl_155 br_155 wl_97 vdd gnd cell_6t
Xbit_r98_c155 bl_155 br_155 wl_98 vdd gnd cell_6t
Xbit_r99_c155 bl_155 br_155 wl_99 vdd gnd cell_6t
Xbit_r100_c155 bl_155 br_155 wl_100 vdd gnd cell_6t
Xbit_r101_c155 bl_155 br_155 wl_101 vdd gnd cell_6t
Xbit_r102_c155 bl_155 br_155 wl_102 vdd gnd cell_6t
Xbit_r103_c155 bl_155 br_155 wl_103 vdd gnd cell_6t
Xbit_r104_c155 bl_155 br_155 wl_104 vdd gnd cell_6t
Xbit_r105_c155 bl_155 br_155 wl_105 vdd gnd cell_6t
Xbit_r106_c155 bl_155 br_155 wl_106 vdd gnd cell_6t
Xbit_r107_c155 bl_155 br_155 wl_107 vdd gnd cell_6t
Xbit_r108_c155 bl_155 br_155 wl_108 vdd gnd cell_6t
Xbit_r109_c155 bl_155 br_155 wl_109 vdd gnd cell_6t
Xbit_r110_c155 bl_155 br_155 wl_110 vdd gnd cell_6t
Xbit_r111_c155 bl_155 br_155 wl_111 vdd gnd cell_6t
Xbit_r112_c155 bl_155 br_155 wl_112 vdd gnd cell_6t
Xbit_r113_c155 bl_155 br_155 wl_113 vdd gnd cell_6t
Xbit_r114_c155 bl_155 br_155 wl_114 vdd gnd cell_6t
Xbit_r115_c155 bl_155 br_155 wl_115 vdd gnd cell_6t
Xbit_r116_c155 bl_155 br_155 wl_116 vdd gnd cell_6t
Xbit_r117_c155 bl_155 br_155 wl_117 vdd gnd cell_6t
Xbit_r118_c155 bl_155 br_155 wl_118 vdd gnd cell_6t
Xbit_r119_c155 bl_155 br_155 wl_119 vdd gnd cell_6t
Xbit_r120_c155 bl_155 br_155 wl_120 vdd gnd cell_6t
Xbit_r121_c155 bl_155 br_155 wl_121 vdd gnd cell_6t
Xbit_r122_c155 bl_155 br_155 wl_122 vdd gnd cell_6t
Xbit_r123_c155 bl_155 br_155 wl_123 vdd gnd cell_6t
Xbit_r124_c155 bl_155 br_155 wl_124 vdd gnd cell_6t
Xbit_r125_c155 bl_155 br_155 wl_125 vdd gnd cell_6t
Xbit_r126_c155 bl_155 br_155 wl_126 vdd gnd cell_6t
Xbit_r127_c155 bl_155 br_155 wl_127 vdd gnd cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd cell_6t
Xbit_r1_c156 bl_156 br_156 wl_1 vdd gnd cell_6t
Xbit_r2_c156 bl_156 br_156 wl_2 vdd gnd cell_6t
Xbit_r3_c156 bl_156 br_156 wl_3 vdd gnd cell_6t
Xbit_r4_c156 bl_156 br_156 wl_4 vdd gnd cell_6t
Xbit_r5_c156 bl_156 br_156 wl_5 vdd gnd cell_6t
Xbit_r6_c156 bl_156 br_156 wl_6 vdd gnd cell_6t
Xbit_r7_c156 bl_156 br_156 wl_7 vdd gnd cell_6t
Xbit_r8_c156 bl_156 br_156 wl_8 vdd gnd cell_6t
Xbit_r9_c156 bl_156 br_156 wl_9 vdd gnd cell_6t
Xbit_r10_c156 bl_156 br_156 wl_10 vdd gnd cell_6t
Xbit_r11_c156 bl_156 br_156 wl_11 vdd gnd cell_6t
Xbit_r12_c156 bl_156 br_156 wl_12 vdd gnd cell_6t
Xbit_r13_c156 bl_156 br_156 wl_13 vdd gnd cell_6t
Xbit_r14_c156 bl_156 br_156 wl_14 vdd gnd cell_6t
Xbit_r15_c156 bl_156 br_156 wl_15 vdd gnd cell_6t
Xbit_r16_c156 bl_156 br_156 wl_16 vdd gnd cell_6t
Xbit_r17_c156 bl_156 br_156 wl_17 vdd gnd cell_6t
Xbit_r18_c156 bl_156 br_156 wl_18 vdd gnd cell_6t
Xbit_r19_c156 bl_156 br_156 wl_19 vdd gnd cell_6t
Xbit_r20_c156 bl_156 br_156 wl_20 vdd gnd cell_6t
Xbit_r21_c156 bl_156 br_156 wl_21 vdd gnd cell_6t
Xbit_r22_c156 bl_156 br_156 wl_22 vdd gnd cell_6t
Xbit_r23_c156 bl_156 br_156 wl_23 vdd gnd cell_6t
Xbit_r24_c156 bl_156 br_156 wl_24 vdd gnd cell_6t
Xbit_r25_c156 bl_156 br_156 wl_25 vdd gnd cell_6t
Xbit_r26_c156 bl_156 br_156 wl_26 vdd gnd cell_6t
Xbit_r27_c156 bl_156 br_156 wl_27 vdd gnd cell_6t
Xbit_r28_c156 bl_156 br_156 wl_28 vdd gnd cell_6t
Xbit_r29_c156 bl_156 br_156 wl_29 vdd gnd cell_6t
Xbit_r30_c156 bl_156 br_156 wl_30 vdd gnd cell_6t
Xbit_r31_c156 bl_156 br_156 wl_31 vdd gnd cell_6t
Xbit_r32_c156 bl_156 br_156 wl_32 vdd gnd cell_6t
Xbit_r33_c156 bl_156 br_156 wl_33 vdd gnd cell_6t
Xbit_r34_c156 bl_156 br_156 wl_34 vdd gnd cell_6t
Xbit_r35_c156 bl_156 br_156 wl_35 vdd gnd cell_6t
Xbit_r36_c156 bl_156 br_156 wl_36 vdd gnd cell_6t
Xbit_r37_c156 bl_156 br_156 wl_37 vdd gnd cell_6t
Xbit_r38_c156 bl_156 br_156 wl_38 vdd gnd cell_6t
Xbit_r39_c156 bl_156 br_156 wl_39 vdd gnd cell_6t
Xbit_r40_c156 bl_156 br_156 wl_40 vdd gnd cell_6t
Xbit_r41_c156 bl_156 br_156 wl_41 vdd gnd cell_6t
Xbit_r42_c156 bl_156 br_156 wl_42 vdd gnd cell_6t
Xbit_r43_c156 bl_156 br_156 wl_43 vdd gnd cell_6t
Xbit_r44_c156 bl_156 br_156 wl_44 vdd gnd cell_6t
Xbit_r45_c156 bl_156 br_156 wl_45 vdd gnd cell_6t
Xbit_r46_c156 bl_156 br_156 wl_46 vdd gnd cell_6t
Xbit_r47_c156 bl_156 br_156 wl_47 vdd gnd cell_6t
Xbit_r48_c156 bl_156 br_156 wl_48 vdd gnd cell_6t
Xbit_r49_c156 bl_156 br_156 wl_49 vdd gnd cell_6t
Xbit_r50_c156 bl_156 br_156 wl_50 vdd gnd cell_6t
Xbit_r51_c156 bl_156 br_156 wl_51 vdd gnd cell_6t
Xbit_r52_c156 bl_156 br_156 wl_52 vdd gnd cell_6t
Xbit_r53_c156 bl_156 br_156 wl_53 vdd gnd cell_6t
Xbit_r54_c156 bl_156 br_156 wl_54 vdd gnd cell_6t
Xbit_r55_c156 bl_156 br_156 wl_55 vdd gnd cell_6t
Xbit_r56_c156 bl_156 br_156 wl_56 vdd gnd cell_6t
Xbit_r57_c156 bl_156 br_156 wl_57 vdd gnd cell_6t
Xbit_r58_c156 bl_156 br_156 wl_58 vdd gnd cell_6t
Xbit_r59_c156 bl_156 br_156 wl_59 vdd gnd cell_6t
Xbit_r60_c156 bl_156 br_156 wl_60 vdd gnd cell_6t
Xbit_r61_c156 bl_156 br_156 wl_61 vdd gnd cell_6t
Xbit_r62_c156 bl_156 br_156 wl_62 vdd gnd cell_6t
Xbit_r63_c156 bl_156 br_156 wl_63 vdd gnd cell_6t
Xbit_r64_c156 bl_156 br_156 wl_64 vdd gnd cell_6t
Xbit_r65_c156 bl_156 br_156 wl_65 vdd gnd cell_6t
Xbit_r66_c156 bl_156 br_156 wl_66 vdd gnd cell_6t
Xbit_r67_c156 bl_156 br_156 wl_67 vdd gnd cell_6t
Xbit_r68_c156 bl_156 br_156 wl_68 vdd gnd cell_6t
Xbit_r69_c156 bl_156 br_156 wl_69 vdd gnd cell_6t
Xbit_r70_c156 bl_156 br_156 wl_70 vdd gnd cell_6t
Xbit_r71_c156 bl_156 br_156 wl_71 vdd gnd cell_6t
Xbit_r72_c156 bl_156 br_156 wl_72 vdd gnd cell_6t
Xbit_r73_c156 bl_156 br_156 wl_73 vdd gnd cell_6t
Xbit_r74_c156 bl_156 br_156 wl_74 vdd gnd cell_6t
Xbit_r75_c156 bl_156 br_156 wl_75 vdd gnd cell_6t
Xbit_r76_c156 bl_156 br_156 wl_76 vdd gnd cell_6t
Xbit_r77_c156 bl_156 br_156 wl_77 vdd gnd cell_6t
Xbit_r78_c156 bl_156 br_156 wl_78 vdd gnd cell_6t
Xbit_r79_c156 bl_156 br_156 wl_79 vdd gnd cell_6t
Xbit_r80_c156 bl_156 br_156 wl_80 vdd gnd cell_6t
Xbit_r81_c156 bl_156 br_156 wl_81 vdd gnd cell_6t
Xbit_r82_c156 bl_156 br_156 wl_82 vdd gnd cell_6t
Xbit_r83_c156 bl_156 br_156 wl_83 vdd gnd cell_6t
Xbit_r84_c156 bl_156 br_156 wl_84 vdd gnd cell_6t
Xbit_r85_c156 bl_156 br_156 wl_85 vdd gnd cell_6t
Xbit_r86_c156 bl_156 br_156 wl_86 vdd gnd cell_6t
Xbit_r87_c156 bl_156 br_156 wl_87 vdd gnd cell_6t
Xbit_r88_c156 bl_156 br_156 wl_88 vdd gnd cell_6t
Xbit_r89_c156 bl_156 br_156 wl_89 vdd gnd cell_6t
Xbit_r90_c156 bl_156 br_156 wl_90 vdd gnd cell_6t
Xbit_r91_c156 bl_156 br_156 wl_91 vdd gnd cell_6t
Xbit_r92_c156 bl_156 br_156 wl_92 vdd gnd cell_6t
Xbit_r93_c156 bl_156 br_156 wl_93 vdd gnd cell_6t
Xbit_r94_c156 bl_156 br_156 wl_94 vdd gnd cell_6t
Xbit_r95_c156 bl_156 br_156 wl_95 vdd gnd cell_6t
Xbit_r96_c156 bl_156 br_156 wl_96 vdd gnd cell_6t
Xbit_r97_c156 bl_156 br_156 wl_97 vdd gnd cell_6t
Xbit_r98_c156 bl_156 br_156 wl_98 vdd gnd cell_6t
Xbit_r99_c156 bl_156 br_156 wl_99 vdd gnd cell_6t
Xbit_r100_c156 bl_156 br_156 wl_100 vdd gnd cell_6t
Xbit_r101_c156 bl_156 br_156 wl_101 vdd gnd cell_6t
Xbit_r102_c156 bl_156 br_156 wl_102 vdd gnd cell_6t
Xbit_r103_c156 bl_156 br_156 wl_103 vdd gnd cell_6t
Xbit_r104_c156 bl_156 br_156 wl_104 vdd gnd cell_6t
Xbit_r105_c156 bl_156 br_156 wl_105 vdd gnd cell_6t
Xbit_r106_c156 bl_156 br_156 wl_106 vdd gnd cell_6t
Xbit_r107_c156 bl_156 br_156 wl_107 vdd gnd cell_6t
Xbit_r108_c156 bl_156 br_156 wl_108 vdd gnd cell_6t
Xbit_r109_c156 bl_156 br_156 wl_109 vdd gnd cell_6t
Xbit_r110_c156 bl_156 br_156 wl_110 vdd gnd cell_6t
Xbit_r111_c156 bl_156 br_156 wl_111 vdd gnd cell_6t
Xbit_r112_c156 bl_156 br_156 wl_112 vdd gnd cell_6t
Xbit_r113_c156 bl_156 br_156 wl_113 vdd gnd cell_6t
Xbit_r114_c156 bl_156 br_156 wl_114 vdd gnd cell_6t
Xbit_r115_c156 bl_156 br_156 wl_115 vdd gnd cell_6t
Xbit_r116_c156 bl_156 br_156 wl_116 vdd gnd cell_6t
Xbit_r117_c156 bl_156 br_156 wl_117 vdd gnd cell_6t
Xbit_r118_c156 bl_156 br_156 wl_118 vdd gnd cell_6t
Xbit_r119_c156 bl_156 br_156 wl_119 vdd gnd cell_6t
Xbit_r120_c156 bl_156 br_156 wl_120 vdd gnd cell_6t
Xbit_r121_c156 bl_156 br_156 wl_121 vdd gnd cell_6t
Xbit_r122_c156 bl_156 br_156 wl_122 vdd gnd cell_6t
Xbit_r123_c156 bl_156 br_156 wl_123 vdd gnd cell_6t
Xbit_r124_c156 bl_156 br_156 wl_124 vdd gnd cell_6t
Xbit_r125_c156 bl_156 br_156 wl_125 vdd gnd cell_6t
Xbit_r126_c156 bl_156 br_156 wl_126 vdd gnd cell_6t
Xbit_r127_c156 bl_156 br_156 wl_127 vdd gnd cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd cell_6t
Xbit_r1_c157 bl_157 br_157 wl_1 vdd gnd cell_6t
Xbit_r2_c157 bl_157 br_157 wl_2 vdd gnd cell_6t
Xbit_r3_c157 bl_157 br_157 wl_3 vdd gnd cell_6t
Xbit_r4_c157 bl_157 br_157 wl_4 vdd gnd cell_6t
Xbit_r5_c157 bl_157 br_157 wl_5 vdd gnd cell_6t
Xbit_r6_c157 bl_157 br_157 wl_6 vdd gnd cell_6t
Xbit_r7_c157 bl_157 br_157 wl_7 vdd gnd cell_6t
Xbit_r8_c157 bl_157 br_157 wl_8 vdd gnd cell_6t
Xbit_r9_c157 bl_157 br_157 wl_9 vdd gnd cell_6t
Xbit_r10_c157 bl_157 br_157 wl_10 vdd gnd cell_6t
Xbit_r11_c157 bl_157 br_157 wl_11 vdd gnd cell_6t
Xbit_r12_c157 bl_157 br_157 wl_12 vdd gnd cell_6t
Xbit_r13_c157 bl_157 br_157 wl_13 vdd gnd cell_6t
Xbit_r14_c157 bl_157 br_157 wl_14 vdd gnd cell_6t
Xbit_r15_c157 bl_157 br_157 wl_15 vdd gnd cell_6t
Xbit_r16_c157 bl_157 br_157 wl_16 vdd gnd cell_6t
Xbit_r17_c157 bl_157 br_157 wl_17 vdd gnd cell_6t
Xbit_r18_c157 bl_157 br_157 wl_18 vdd gnd cell_6t
Xbit_r19_c157 bl_157 br_157 wl_19 vdd gnd cell_6t
Xbit_r20_c157 bl_157 br_157 wl_20 vdd gnd cell_6t
Xbit_r21_c157 bl_157 br_157 wl_21 vdd gnd cell_6t
Xbit_r22_c157 bl_157 br_157 wl_22 vdd gnd cell_6t
Xbit_r23_c157 bl_157 br_157 wl_23 vdd gnd cell_6t
Xbit_r24_c157 bl_157 br_157 wl_24 vdd gnd cell_6t
Xbit_r25_c157 bl_157 br_157 wl_25 vdd gnd cell_6t
Xbit_r26_c157 bl_157 br_157 wl_26 vdd gnd cell_6t
Xbit_r27_c157 bl_157 br_157 wl_27 vdd gnd cell_6t
Xbit_r28_c157 bl_157 br_157 wl_28 vdd gnd cell_6t
Xbit_r29_c157 bl_157 br_157 wl_29 vdd gnd cell_6t
Xbit_r30_c157 bl_157 br_157 wl_30 vdd gnd cell_6t
Xbit_r31_c157 bl_157 br_157 wl_31 vdd gnd cell_6t
Xbit_r32_c157 bl_157 br_157 wl_32 vdd gnd cell_6t
Xbit_r33_c157 bl_157 br_157 wl_33 vdd gnd cell_6t
Xbit_r34_c157 bl_157 br_157 wl_34 vdd gnd cell_6t
Xbit_r35_c157 bl_157 br_157 wl_35 vdd gnd cell_6t
Xbit_r36_c157 bl_157 br_157 wl_36 vdd gnd cell_6t
Xbit_r37_c157 bl_157 br_157 wl_37 vdd gnd cell_6t
Xbit_r38_c157 bl_157 br_157 wl_38 vdd gnd cell_6t
Xbit_r39_c157 bl_157 br_157 wl_39 vdd gnd cell_6t
Xbit_r40_c157 bl_157 br_157 wl_40 vdd gnd cell_6t
Xbit_r41_c157 bl_157 br_157 wl_41 vdd gnd cell_6t
Xbit_r42_c157 bl_157 br_157 wl_42 vdd gnd cell_6t
Xbit_r43_c157 bl_157 br_157 wl_43 vdd gnd cell_6t
Xbit_r44_c157 bl_157 br_157 wl_44 vdd gnd cell_6t
Xbit_r45_c157 bl_157 br_157 wl_45 vdd gnd cell_6t
Xbit_r46_c157 bl_157 br_157 wl_46 vdd gnd cell_6t
Xbit_r47_c157 bl_157 br_157 wl_47 vdd gnd cell_6t
Xbit_r48_c157 bl_157 br_157 wl_48 vdd gnd cell_6t
Xbit_r49_c157 bl_157 br_157 wl_49 vdd gnd cell_6t
Xbit_r50_c157 bl_157 br_157 wl_50 vdd gnd cell_6t
Xbit_r51_c157 bl_157 br_157 wl_51 vdd gnd cell_6t
Xbit_r52_c157 bl_157 br_157 wl_52 vdd gnd cell_6t
Xbit_r53_c157 bl_157 br_157 wl_53 vdd gnd cell_6t
Xbit_r54_c157 bl_157 br_157 wl_54 vdd gnd cell_6t
Xbit_r55_c157 bl_157 br_157 wl_55 vdd gnd cell_6t
Xbit_r56_c157 bl_157 br_157 wl_56 vdd gnd cell_6t
Xbit_r57_c157 bl_157 br_157 wl_57 vdd gnd cell_6t
Xbit_r58_c157 bl_157 br_157 wl_58 vdd gnd cell_6t
Xbit_r59_c157 bl_157 br_157 wl_59 vdd gnd cell_6t
Xbit_r60_c157 bl_157 br_157 wl_60 vdd gnd cell_6t
Xbit_r61_c157 bl_157 br_157 wl_61 vdd gnd cell_6t
Xbit_r62_c157 bl_157 br_157 wl_62 vdd gnd cell_6t
Xbit_r63_c157 bl_157 br_157 wl_63 vdd gnd cell_6t
Xbit_r64_c157 bl_157 br_157 wl_64 vdd gnd cell_6t
Xbit_r65_c157 bl_157 br_157 wl_65 vdd gnd cell_6t
Xbit_r66_c157 bl_157 br_157 wl_66 vdd gnd cell_6t
Xbit_r67_c157 bl_157 br_157 wl_67 vdd gnd cell_6t
Xbit_r68_c157 bl_157 br_157 wl_68 vdd gnd cell_6t
Xbit_r69_c157 bl_157 br_157 wl_69 vdd gnd cell_6t
Xbit_r70_c157 bl_157 br_157 wl_70 vdd gnd cell_6t
Xbit_r71_c157 bl_157 br_157 wl_71 vdd gnd cell_6t
Xbit_r72_c157 bl_157 br_157 wl_72 vdd gnd cell_6t
Xbit_r73_c157 bl_157 br_157 wl_73 vdd gnd cell_6t
Xbit_r74_c157 bl_157 br_157 wl_74 vdd gnd cell_6t
Xbit_r75_c157 bl_157 br_157 wl_75 vdd gnd cell_6t
Xbit_r76_c157 bl_157 br_157 wl_76 vdd gnd cell_6t
Xbit_r77_c157 bl_157 br_157 wl_77 vdd gnd cell_6t
Xbit_r78_c157 bl_157 br_157 wl_78 vdd gnd cell_6t
Xbit_r79_c157 bl_157 br_157 wl_79 vdd gnd cell_6t
Xbit_r80_c157 bl_157 br_157 wl_80 vdd gnd cell_6t
Xbit_r81_c157 bl_157 br_157 wl_81 vdd gnd cell_6t
Xbit_r82_c157 bl_157 br_157 wl_82 vdd gnd cell_6t
Xbit_r83_c157 bl_157 br_157 wl_83 vdd gnd cell_6t
Xbit_r84_c157 bl_157 br_157 wl_84 vdd gnd cell_6t
Xbit_r85_c157 bl_157 br_157 wl_85 vdd gnd cell_6t
Xbit_r86_c157 bl_157 br_157 wl_86 vdd gnd cell_6t
Xbit_r87_c157 bl_157 br_157 wl_87 vdd gnd cell_6t
Xbit_r88_c157 bl_157 br_157 wl_88 vdd gnd cell_6t
Xbit_r89_c157 bl_157 br_157 wl_89 vdd gnd cell_6t
Xbit_r90_c157 bl_157 br_157 wl_90 vdd gnd cell_6t
Xbit_r91_c157 bl_157 br_157 wl_91 vdd gnd cell_6t
Xbit_r92_c157 bl_157 br_157 wl_92 vdd gnd cell_6t
Xbit_r93_c157 bl_157 br_157 wl_93 vdd gnd cell_6t
Xbit_r94_c157 bl_157 br_157 wl_94 vdd gnd cell_6t
Xbit_r95_c157 bl_157 br_157 wl_95 vdd gnd cell_6t
Xbit_r96_c157 bl_157 br_157 wl_96 vdd gnd cell_6t
Xbit_r97_c157 bl_157 br_157 wl_97 vdd gnd cell_6t
Xbit_r98_c157 bl_157 br_157 wl_98 vdd gnd cell_6t
Xbit_r99_c157 bl_157 br_157 wl_99 vdd gnd cell_6t
Xbit_r100_c157 bl_157 br_157 wl_100 vdd gnd cell_6t
Xbit_r101_c157 bl_157 br_157 wl_101 vdd gnd cell_6t
Xbit_r102_c157 bl_157 br_157 wl_102 vdd gnd cell_6t
Xbit_r103_c157 bl_157 br_157 wl_103 vdd gnd cell_6t
Xbit_r104_c157 bl_157 br_157 wl_104 vdd gnd cell_6t
Xbit_r105_c157 bl_157 br_157 wl_105 vdd gnd cell_6t
Xbit_r106_c157 bl_157 br_157 wl_106 vdd gnd cell_6t
Xbit_r107_c157 bl_157 br_157 wl_107 vdd gnd cell_6t
Xbit_r108_c157 bl_157 br_157 wl_108 vdd gnd cell_6t
Xbit_r109_c157 bl_157 br_157 wl_109 vdd gnd cell_6t
Xbit_r110_c157 bl_157 br_157 wl_110 vdd gnd cell_6t
Xbit_r111_c157 bl_157 br_157 wl_111 vdd gnd cell_6t
Xbit_r112_c157 bl_157 br_157 wl_112 vdd gnd cell_6t
Xbit_r113_c157 bl_157 br_157 wl_113 vdd gnd cell_6t
Xbit_r114_c157 bl_157 br_157 wl_114 vdd gnd cell_6t
Xbit_r115_c157 bl_157 br_157 wl_115 vdd gnd cell_6t
Xbit_r116_c157 bl_157 br_157 wl_116 vdd gnd cell_6t
Xbit_r117_c157 bl_157 br_157 wl_117 vdd gnd cell_6t
Xbit_r118_c157 bl_157 br_157 wl_118 vdd gnd cell_6t
Xbit_r119_c157 bl_157 br_157 wl_119 vdd gnd cell_6t
Xbit_r120_c157 bl_157 br_157 wl_120 vdd gnd cell_6t
Xbit_r121_c157 bl_157 br_157 wl_121 vdd gnd cell_6t
Xbit_r122_c157 bl_157 br_157 wl_122 vdd gnd cell_6t
Xbit_r123_c157 bl_157 br_157 wl_123 vdd gnd cell_6t
Xbit_r124_c157 bl_157 br_157 wl_124 vdd gnd cell_6t
Xbit_r125_c157 bl_157 br_157 wl_125 vdd gnd cell_6t
Xbit_r126_c157 bl_157 br_157 wl_126 vdd gnd cell_6t
Xbit_r127_c157 bl_157 br_157 wl_127 vdd gnd cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd cell_6t
Xbit_r1_c158 bl_158 br_158 wl_1 vdd gnd cell_6t
Xbit_r2_c158 bl_158 br_158 wl_2 vdd gnd cell_6t
Xbit_r3_c158 bl_158 br_158 wl_3 vdd gnd cell_6t
Xbit_r4_c158 bl_158 br_158 wl_4 vdd gnd cell_6t
Xbit_r5_c158 bl_158 br_158 wl_5 vdd gnd cell_6t
Xbit_r6_c158 bl_158 br_158 wl_6 vdd gnd cell_6t
Xbit_r7_c158 bl_158 br_158 wl_7 vdd gnd cell_6t
Xbit_r8_c158 bl_158 br_158 wl_8 vdd gnd cell_6t
Xbit_r9_c158 bl_158 br_158 wl_9 vdd gnd cell_6t
Xbit_r10_c158 bl_158 br_158 wl_10 vdd gnd cell_6t
Xbit_r11_c158 bl_158 br_158 wl_11 vdd gnd cell_6t
Xbit_r12_c158 bl_158 br_158 wl_12 vdd gnd cell_6t
Xbit_r13_c158 bl_158 br_158 wl_13 vdd gnd cell_6t
Xbit_r14_c158 bl_158 br_158 wl_14 vdd gnd cell_6t
Xbit_r15_c158 bl_158 br_158 wl_15 vdd gnd cell_6t
Xbit_r16_c158 bl_158 br_158 wl_16 vdd gnd cell_6t
Xbit_r17_c158 bl_158 br_158 wl_17 vdd gnd cell_6t
Xbit_r18_c158 bl_158 br_158 wl_18 vdd gnd cell_6t
Xbit_r19_c158 bl_158 br_158 wl_19 vdd gnd cell_6t
Xbit_r20_c158 bl_158 br_158 wl_20 vdd gnd cell_6t
Xbit_r21_c158 bl_158 br_158 wl_21 vdd gnd cell_6t
Xbit_r22_c158 bl_158 br_158 wl_22 vdd gnd cell_6t
Xbit_r23_c158 bl_158 br_158 wl_23 vdd gnd cell_6t
Xbit_r24_c158 bl_158 br_158 wl_24 vdd gnd cell_6t
Xbit_r25_c158 bl_158 br_158 wl_25 vdd gnd cell_6t
Xbit_r26_c158 bl_158 br_158 wl_26 vdd gnd cell_6t
Xbit_r27_c158 bl_158 br_158 wl_27 vdd gnd cell_6t
Xbit_r28_c158 bl_158 br_158 wl_28 vdd gnd cell_6t
Xbit_r29_c158 bl_158 br_158 wl_29 vdd gnd cell_6t
Xbit_r30_c158 bl_158 br_158 wl_30 vdd gnd cell_6t
Xbit_r31_c158 bl_158 br_158 wl_31 vdd gnd cell_6t
Xbit_r32_c158 bl_158 br_158 wl_32 vdd gnd cell_6t
Xbit_r33_c158 bl_158 br_158 wl_33 vdd gnd cell_6t
Xbit_r34_c158 bl_158 br_158 wl_34 vdd gnd cell_6t
Xbit_r35_c158 bl_158 br_158 wl_35 vdd gnd cell_6t
Xbit_r36_c158 bl_158 br_158 wl_36 vdd gnd cell_6t
Xbit_r37_c158 bl_158 br_158 wl_37 vdd gnd cell_6t
Xbit_r38_c158 bl_158 br_158 wl_38 vdd gnd cell_6t
Xbit_r39_c158 bl_158 br_158 wl_39 vdd gnd cell_6t
Xbit_r40_c158 bl_158 br_158 wl_40 vdd gnd cell_6t
Xbit_r41_c158 bl_158 br_158 wl_41 vdd gnd cell_6t
Xbit_r42_c158 bl_158 br_158 wl_42 vdd gnd cell_6t
Xbit_r43_c158 bl_158 br_158 wl_43 vdd gnd cell_6t
Xbit_r44_c158 bl_158 br_158 wl_44 vdd gnd cell_6t
Xbit_r45_c158 bl_158 br_158 wl_45 vdd gnd cell_6t
Xbit_r46_c158 bl_158 br_158 wl_46 vdd gnd cell_6t
Xbit_r47_c158 bl_158 br_158 wl_47 vdd gnd cell_6t
Xbit_r48_c158 bl_158 br_158 wl_48 vdd gnd cell_6t
Xbit_r49_c158 bl_158 br_158 wl_49 vdd gnd cell_6t
Xbit_r50_c158 bl_158 br_158 wl_50 vdd gnd cell_6t
Xbit_r51_c158 bl_158 br_158 wl_51 vdd gnd cell_6t
Xbit_r52_c158 bl_158 br_158 wl_52 vdd gnd cell_6t
Xbit_r53_c158 bl_158 br_158 wl_53 vdd gnd cell_6t
Xbit_r54_c158 bl_158 br_158 wl_54 vdd gnd cell_6t
Xbit_r55_c158 bl_158 br_158 wl_55 vdd gnd cell_6t
Xbit_r56_c158 bl_158 br_158 wl_56 vdd gnd cell_6t
Xbit_r57_c158 bl_158 br_158 wl_57 vdd gnd cell_6t
Xbit_r58_c158 bl_158 br_158 wl_58 vdd gnd cell_6t
Xbit_r59_c158 bl_158 br_158 wl_59 vdd gnd cell_6t
Xbit_r60_c158 bl_158 br_158 wl_60 vdd gnd cell_6t
Xbit_r61_c158 bl_158 br_158 wl_61 vdd gnd cell_6t
Xbit_r62_c158 bl_158 br_158 wl_62 vdd gnd cell_6t
Xbit_r63_c158 bl_158 br_158 wl_63 vdd gnd cell_6t
Xbit_r64_c158 bl_158 br_158 wl_64 vdd gnd cell_6t
Xbit_r65_c158 bl_158 br_158 wl_65 vdd gnd cell_6t
Xbit_r66_c158 bl_158 br_158 wl_66 vdd gnd cell_6t
Xbit_r67_c158 bl_158 br_158 wl_67 vdd gnd cell_6t
Xbit_r68_c158 bl_158 br_158 wl_68 vdd gnd cell_6t
Xbit_r69_c158 bl_158 br_158 wl_69 vdd gnd cell_6t
Xbit_r70_c158 bl_158 br_158 wl_70 vdd gnd cell_6t
Xbit_r71_c158 bl_158 br_158 wl_71 vdd gnd cell_6t
Xbit_r72_c158 bl_158 br_158 wl_72 vdd gnd cell_6t
Xbit_r73_c158 bl_158 br_158 wl_73 vdd gnd cell_6t
Xbit_r74_c158 bl_158 br_158 wl_74 vdd gnd cell_6t
Xbit_r75_c158 bl_158 br_158 wl_75 vdd gnd cell_6t
Xbit_r76_c158 bl_158 br_158 wl_76 vdd gnd cell_6t
Xbit_r77_c158 bl_158 br_158 wl_77 vdd gnd cell_6t
Xbit_r78_c158 bl_158 br_158 wl_78 vdd gnd cell_6t
Xbit_r79_c158 bl_158 br_158 wl_79 vdd gnd cell_6t
Xbit_r80_c158 bl_158 br_158 wl_80 vdd gnd cell_6t
Xbit_r81_c158 bl_158 br_158 wl_81 vdd gnd cell_6t
Xbit_r82_c158 bl_158 br_158 wl_82 vdd gnd cell_6t
Xbit_r83_c158 bl_158 br_158 wl_83 vdd gnd cell_6t
Xbit_r84_c158 bl_158 br_158 wl_84 vdd gnd cell_6t
Xbit_r85_c158 bl_158 br_158 wl_85 vdd gnd cell_6t
Xbit_r86_c158 bl_158 br_158 wl_86 vdd gnd cell_6t
Xbit_r87_c158 bl_158 br_158 wl_87 vdd gnd cell_6t
Xbit_r88_c158 bl_158 br_158 wl_88 vdd gnd cell_6t
Xbit_r89_c158 bl_158 br_158 wl_89 vdd gnd cell_6t
Xbit_r90_c158 bl_158 br_158 wl_90 vdd gnd cell_6t
Xbit_r91_c158 bl_158 br_158 wl_91 vdd gnd cell_6t
Xbit_r92_c158 bl_158 br_158 wl_92 vdd gnd cell_6t
Xbit_r93_c158 bl_158 br_158 wl_93 vdd gnd cell_6t
Xbit_r94_c158 bl_158 br_158 wl_94 vdd gnd cell_6t
Xbit_r95_c158 bl_158 br_158 wl_95 vdd gnd cell_6t
Xbit_r96_c158 bl_158 br_158 wl_96 vdd gnd cell_6t
Xbit_r97_c158 bl_158 br_158 wl_97 vdd gnd cell_6t
Xbit_r98_c158 bl_158 br_158 wl_98 vdd gnd cell_6t
Xbit_r99_c158 bl_158 br_158 wl_99 vdd gnd cell_6t
Xbit_r100_c158 bl_158 br_158 wl_100 vdd gnd cell_6t
Xbit_r101_c158 bl_158 br_158 wl_101 vdd gnd cell_6t
Xbit_r102_c158 bl_158 br_158 wl_102 vdd gnd cell_6t
Xbit_r103_c158 bl_158 br_158 wl_103 vdd gnd cell_6t
Xbit_r104_c158 bl_158 br_158 wl_104 vdd gnd cell_6t
Xbit_r105_c158 bl_158 br_158 wl_105 vdd gnd cell_6t
Xbit_r106_c158 bl_158 br_158 wl_106 vdd gnd cell_6t
Xbit_r107_c158 bl_158 br_158 wl_107 vdd gnd cell_6t
Xbit_r108_c158 bl_158 br_158 wl_108 vdd gnd cell_6t
Xbit_r109_c158 bl_158 br_158 wl_109 vdd gnd cell_6t
Xbit_r110_c158 bl_158 br_158 wl_110 vdd gnd cell_6t
Xbit_r111_c158 bl_158 br_158 wl_111 vdd gnd cell_6t
Xbit_r112_c158 bl_158 br_158 wl_112 vdd gnd cell_6t
Xbit_r113_c158 bl_158 br_158 wl_113 vdd gnd cell_6t
Xbit_r114_c158 bl_158 br_158 wl_114 vdd gnd cell_6t
Xbit_r115_c158 bl_158 br_158 wl_115 vdd gnd cell_6t
Xbit_r116_c158 bl_158 br_158 wl_116 vdd gnd cell_6t
Xbit_r117_c158 bl_158 br_158 wl_117 vdd gnd cell_6t
Xbit_r118_c158 bl_158 br_158 wl_118 vdd gnd cell_6t
Xbit_r119_c158 bl_158 br_158 wl_119 vdd gnd cell_6t
Xbit_r120_c158 bl_158 br_158 wl_120 vdd gnd cell_6t
Xbit_r121_c158 bl_158 br_158 wl_121 vdd gnd cell_6t
Xbit_r122_c158 bl_158 br_158 wl_122 vdd gnd cell_6t
Xbit_r123_c158 bl_158 br_158 wl_123 vdd gnd cell_6t
Xbit_r124_c158 bl_158 br_158 wl_124 vdd gnd cell_6t
Xbit_r125_c158 bl_158 br_158 wl_125 vdd gnd cell_6t
Xbit_r126_c158 bl_158 br_158 wl_126 vdd gnd cell_6t
Xbit_r127_c158 bl_158 br_158 wl_127 vdd gnd cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd cell_6t
Xbit_r1_c159 bl_159 br_159 wl_1 vdd gnd cell_6t
Xbit_r2_c159 bl_159 br_159 wl_2 vdd gnd cell_6t
Xbit_r3_c159 bl_159 br_159 wl_3 vdd gnd cell_6t
Xbit_r4_c159 bl_159 br_159 wl_4 vdd gnd cell_6t
Xbit_r5_c159 bl_159 br_159 wl_5 vdd gnd cell_6t
Xbit_r6_c159 bl_159 br_159 wl_6 vdd gnd cell_6t
Xbit_r7_c159 bl_159 br_159 wl_7 vdd gnd cell_6t
Xbit_r8_c159 bl_159 br_159 wl_8 vdd gnd cell_6t
Xbit_r9_c159 bl_159 br_159 wl_9 vdd gnd cell_6t
Xbit_r10_c159 bl_159 br_159 wl_10 vdd gnd cell_6t
Xbit_r11_c159 bl_159 br_159 wl_11 vdd gnd cell_6t
Xbit_r12_c159 bl_159 br_159 wl_12 vdd gnd cell_6t
Xbit_r13_c159 bl_159 br_159 wl_13 vdd gnd cell_6t
Xbit_r14_c159 bl_159 br_159 wl_14 vdd gnd cell_6t
Xbit_r15_c159 bl_159 br_159 wl_15 vdd gnd cell_6t
Xbit_r16_c159 bl_159 br_159 wl_16 vdd gnd cell_6t
Xbit_r17_c159 bl_159 br_159 wl_17 vdd gnd cell_6t
Xbit_r18_c159 bl_159 br_159 wl_18 vdd gnd cell_6t
Xbit_r19_c159 bl_159 br_159 wl_19 vdd gnd cell_6t
Xbit_r20_c159 bl_159 br_159 wl_20 vdd gnd cell_6t
Xbit_r21_c159 bl_159 br_159 wl_21 vdd gnd cell_6t
Xbit_r22_c159 bl_159 br_159 wl_22 vdd gnd cell_6t
Xbit_r23_c159 bl_159 br_159 wl_23 vdd gnd cell_6t
Xbit_r24_c159 bl_159 br_159 wl_24 vdd gnd cell_6t
Xbit_r25_c159 bl_159 br_159 wl_25 vdd gnd cell_6t
Xbit_r26_c159 bl_159 br_159 wl_26 vdd gnd cell_6t
Xbit_r27_c159 bl_159 br_159 wl_27 vdd gnd cell_6t
Xbit_r28_c159 bl_159 br_159 wl_28 vdd gnd cell_6t
Xbit_r29_c159 bl_159 br_159 wl_29 vdd gnd cell_6t
Xbit_r30_c159 bl_159 br_159 wl_30 vdd gnd cell_6t
Xbit_r31_c159 bl_159 br_159 wl_31 vdd gnd cell_6t
Xbit_r32_c159 bl_159 br_159 wl_32 vdd gnd cell_6t
Xbit_r33_c159 bl_159 br_159 wl_33 vdd gnd cell_6t
Xbit_r34_c159 bl_159 br_159 wl_34 vdd gnd cell_6t
Xbit_r35_c159 bl_159 br_159 wl_35 vdd gnd cell_6t
Xbit_r36_c159 bl_159 br_159 wl_36 vdd gnd cell_6t
Xbit_r37_c159 bl_159 br_159 wl_37 vdd gnd cell_6t
Xbit_r38_c159 bl_159 br_159 wl_38 vdd gnd cell_6t
Xbit_r39_c159 bl_159 br_159 wl_39 vdd gnd cell_6t
Xbit_r40_c159 bl_159 br_159 wl_40 vdd gnd cell_6t
Xbit_r41_c159 bl_159 br_159 wl_41 vdd gnd cell_6t
Xbit_r42_c159 bl_159 br_159 wl_42 vdd gnd cell_6t
Xbit_r43_c159 bl_159 br_159 wl_43 vdd gnd cell_6t
Xbit_r44_c159 bl_159 br_159 wl_44 vdd gnd cell_6t
Xbit_r45_c159 bl_159 br_159 wl_45 vdd gnd cell_6t
Xbit_r46_c159 bl_159 br_159 wl_46 vdd gnd cell_6t
Xbit_r47_c159 bl_159 br_159 wl_47 vdd gnd cell_6t
Xbit_r48_c159 bl_159 br_159 wl_48 vdd gnd cell_6t
Xbit_r49_c159 bl_159 br_159 wl_49 vdd gnd cell_6t
Xbit_r50_c159 bl_159 br_159 wl_50 vdd gnd cell_6t
Xbit_r51_c159 bl_159 br_159 wl_51 vdd gnd cell_6t
Xbit_r52_c159 bl_159 br_159 wl_52 vdd gnd cell_6t
Xbit_r53_c159 bl_159 br_159 wl_53 vdd gnd cell_6t
Xbit_r54_c159 bl_159 br_159 wl_54 vdd gnd cell_6t
Xbit_r55_c159 bl_159 br_159 wl_55 vdd gnd cell_6t
Xbit_r56_c159 bl_159 br_159 wl_56 vdd gnd cell_6t
Xbit_r57_c159 bl_159 br_159 wl_57 vdd gnd cell_6t
Xbit_r58_c159 bl_159 br_159 wl_58 vdd gnd cell_6t
Xbit_r59_c159 bl_159 br_159 wl_59 vdd gnd cell_6t
Xbit_r60_c159 bl_159 br_159 wl_60 vdd gnd cell_6t
Xbit_r61_c159 bl_159 br_159 wl_61 vdd gnd cell_6t
Xbit_r62_c159 bl_159 br_159 wl_62 vdd gnd cell_6t
Xbit_r63_c159 bl_159 br_159 wl_63 vdd gnd cell_6t
Xbit_r64_c159 bl_159 br_159 wl_64 vdd gnd cell_6t
Xbit_r65_c159 bl_159 br_159 wl_65 vdd gnd cell_6t
Xbit_r66_c159 bl_159 br_159 wl_66 vdd gnd cell_6t
Xbit_r67_c159 bl_159 br_159 wl_67 vdd gnd cell_6t
Xbit_r68_c159 bl_159 br_159 wl_68 vdd gnd cell_6t
Xbit_r69_c159 bl_159 br_159 wl_69 vdd gnd cell_6t
Xbit_r70_c159 bl_159 br_159 wl_70 vdd gnd cell_6t
Xbit_r71_c159 bl_159 br_159 wl_71 vdd gnd cell_6t
Xbit_r72_c159 bl_159 br_159 wl_72 vdd gnd cell_6t
Xbit_r73_c159 bl_159 br_159 wl_73 vdd gnd cell_6t
Xbit_r74_c159 bl_159 br_159 wl_74 vdd gnd cell_6t
Xbit_r75_c159 bl_159 br_159 wl_75 vdd gnd cell_6t
Xbit_r76_c159 bl_159 br_159 wl_76 vdd gnd cell_6t
Xbit_r77_c159 bl_159 br_159 wl_77 vdd gnd cell_6t
Xbit_r78_c159 bl_159 br_159 wl_78 vdd gnd cell_6t
Xbit_r79_c159 bl_159 br_159 wl_79 vdd gnd cell_6t
Xbit_r80_c159 bl_159 br_159 wl_80 vdd gnd cell_6t
Xbit_r81_c159 bl_159 br_159 wl_81 vdd gnd cell_6t
Xbit_r82_c159 bl_159 br_159 wl_82 vdd gnd cell_6t
Xbit_r83_c159 bl_159 br_159 wl_83 vdd gnd cell_6t
Xbit_r84_c159 bl_159 br_159 wl_84 vdd gnd cell_6t
Xbit_r85_c159 bl_159 br_159 wl_85 vdd gnd cell_6t
Xbit_r86_c159 bl_159 br_159 wl_86 vdd gnd cell_6t
Xbit_r87_c159 bl_159 br_159 wl_87 vdd gnd cell_6t
Xbit_r88_c159 bl_159 br_159 wl_88 vdd gnd cell_6t
Xbit_r89_c159 bl_159 br_159 wl_89 vdd gnd cell_6t
Xbit_r90_c159 bl_159 br_159 wl_90 vdd gnd cell_6t
Xbit_r91_c159 bl_159 br_159 wl_91 vdd gnd cell_6t
Xbit_r92_c159 bl_159 br_159 wl_92 vdd gnd cell_6t
Xbit_r93_c159 bl_159 br_159 wl_93 vdd gnd cell_6t
Xbit_r94_c159 bl_159 br_159 wl_94 vdd gnd cell_6t
Xbit_r95_c159 bl_159 br_159 wl_95 vdd gnd cell_6t
Xbit_r96_c159 bl_159 br_159 wl_96 vdd gnd cell_6t
Xbit_r97_c159 bl_159 br_159 wl_97 vdd gnd cell_6t
Xbit_r98_c159 bl_159 br_159 wl_98 vdd gnd cell_6t
Xbit_r99_c159 bl_159 br_159 wl_99 vdd gnd cell_6t
Xbit_r100_c159 bl_159 br_159 wl_100 vdd gnd cell_6t
Xbit_r101_c159 bl_159 br_159 wl_101 vdd gnd cell_6t
Xbit_r102_c159 bl_159 br_159 wl_102 vdd gnd cell_6t
Xbit_r103_c159 bl_159 br_159 wl_103 vdd gnd cell_6t
Xbit_r104_c159 bl_159 br_159 wl_104 vdd gnd cell_6t
Xbit_r105_c159 bl_159 br_159 wl_105 vdd gnd cell_6t
Xbit_r106_c159 bl_159 br_159 wl_106 vdd gnd cell_6t
Xbit_r107_c159 bl_159 br_159 wl_107 vdd gnd cell_6t
Xbit_r108_c159 bl_159 br_159 wl_108 vdd gnd cell_6t
Xbit_r109_c159 bl_159 br_159 wl_109 vdd gnd cell_6t
Xbit_r110_c159 bl_159 br_159 wl_110 vdd gnd cell_6t
Xbit_r111_c159 bl_159 br_159 wl_111 vdd gnd cell_6t
Xbit_r112_c159 bl_159 br_159 wl_112 vdd gnd cell_6t
Xbit_r113_c159 bl_159 br_159 wl_113 vdd gnd cell_6t
Xbit_r114_c159 bl_159 br_159 wl_114 vdd gnd cell_6t
Xbit_r115_c159 bl_159 br_159 wl_115 vdd gnd cell_6t
Xbit_r116_c159 bl_159 br_159 wl_116 vdd gnd cell_6t
Xbit_r117_c159 bl_159 br_159 wl_117 vdd gnd cell_6t
Xbit_r118_c159 bl_159 br_159 wl_118 vdd gnd cell_6t
Xbit_r119_c159 bl_159 br_159 wl_119 vdd gnd cell_6t
Xbit_r120_c159 bl_159 br_159 wl_120 vdd gnd cell_6t
Xbit_r121_c159 bl_159 br_159 wl_121 vdd gnd cell_6t
Xbit_r122_c159 bl_159 br_159 wl_122 vdd gnd cell_6t
Xbit_r123_c159 bl_159 br_159 wl_123 vdd gnd cell_6t
Xbit_r124_c159 bl_159 br_159 wl_124 vdd gnd cell_6t
Xbit_r125_c159 bl_159 br_159 wl_125 vdd gnd cell_6t
Xbit_r126_c159 bl_159 br_159 wl_126 vdd gnd cell_6t
Xbit_r127_c159 bl_159 br_159 wl_127 vdd gnd cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd cell_6t
Xbit_r1_c160 bl_160 br_160 wl_1 vdd gnd cell_6t
Xbit_r2_c160 bl_160 br_160 wl_2 vdd gnd cell_6t
Xbit_r3_c160 bl_160 br_160 wl_3 vdd gnd cell_6t
Xbit_r4_c160 bl_160 br_160 wl_4 vdd gnd cell_6t
Xbit_r5_c160 bl_160 br_160 wl_5 vdd gnd cell_6t
Xbit_r6_c160 bl_160 br_160 wl_6 vdd gnd cell_6t
Xbit_r7_c160 bl_160 br_160 wl_7 vdd gnd cell_6t
Xbit_r8_c160 bl_160 br_160 wl_8 vdd gnd cell_6t
Xbit_r9_c160 bl_160 br_160 wl_9 vdd gnd cell_6t
Xbit_r10_c160 bl_160 br_160 wl_10 vdd gnd cell_6t
Xbit_r11_c160 bl_160 br_160 wl_11 vdd gnd cell_6t
Xbit_r12_c160 bl_160 br_160 wl_12 vdd gnd cell_6t
Xbit_r13_c160 bl_160 br_160 wl_13 vdd gnd cell_6t
Xbit_r14_c160 bl_160 br_160 wl_14 vdd gnd cell_6t
Xbit_r15_c160 bl_160 br_160 wl_15 vdd gnd cell_6t
Xbit_r16_c160 bl_160 br_160 wl_16 vdd gnd cell_6t
Xbit_r17_c160 bl_160 br_160 wl_17 vdd gnd cell_6t
Xbit_r18_c160 bl_160 br_160 wl_18 vdd gnd cell_6t
Xbit_r19_c160 bl_160 br_160 wl_19 vdd gnd cell_6t
Xbit_r20_c160 bl_160 br_160 wl_20 vdd gnd cell_6t
Xbit_r21_c160 bl_160 br_160 wl_21 vdd gnd cell_6t
Xbit_r22_c160 bl_160 br_160 wl_22 vdd gnd cell_6t
Xbit_r23_c160 bl_160 br_160 wl_23 vdd gnd cell_6t
Xbit_r24_c160 bl_160 br_160 wl_24 vdd gnd cell_6t
Xbit_r25_c160 bl_160 br_160 wl_25 vdd gnd cell_6t
Xbit_r26_c160 bl_160 br_160 wl_26 vdd gnd cell_6t
Xbit_r27_c160 bl_160 br_160 wl_27 vdd gnd cell_6t
Xbit_r28_c160 bl_160 br_160 wl_28 vdd gnd cell_6t
Xbit_r29_c160 bl_160 br_160 wl_29 vdd gnd cell_6t
Xbit_r30_c160 bl_160 br_160 wl_30 vdd gnd cell_6t
Xbit_r31_c160 bl_160 br_160 wl_31 vdd gnd cell_6t
Xbit_r32_c160 bl_160 br_160 wl_32 vdd gnd cell_6t
Xbit_r33_c160 bl_160 br_160 wl_33 vdd gnd cell_6t
Xbit_r34_c160 bl_160 br_160 wl_34 vdd gnd cell_6t
Xbit_r35_c160 bl_160 br_160 wl_35 vdd gnd cell_6t
Xbit_r36_c160 bl_160 br_160 wl_36 vdd gnd cell_6t
Xbit_r37_c160 bl_160 br_160 wl_37 vdd gnd cell_6t
Xbit_r38_c160 bl_160 br_160 wl_38 vdd gnd cell_6t
Xbit_r39_c160 bl_160 br_160 wl_39 vdd gnd cell_6t
Xbit_r40_c160 bl_160 br_160 wl_40 vdd gnd cell_6t
Xbit_r41_c160 bl_160 br_160 wl_41 vdd gnd cell_6t
Xbit_r42_c160 bl_160 br_160 wl_42 vdd gnd cell_6t
Xbit_r43_c160 bl_160 br_160 wl_43 vdd gnd cell_6t
Xbit_r44_c160 bl_160 br_160 wl_44 vdd gnd cell_6t
Xbit_r45_c160 bl_160 br_160 wl_45 vdd gnd cell_6t
Xbit_r46_c160 bl_160 br_160 wl_46 vdd gnd cell_6t
Xbit_r47_c160 bl_160 br_160 wl_47 vdd gnd cell_6t
Xbit_r48_c160 bl_160 br_160 wl_48 vdd gnd cell_6t
Xbit_r49_c160 bl_160 br_160 wl_49 vdd gnd cell_6t
Xbit_r50_c160 bl_160 br_160 wl_50 vdd gnd cell_6t
Xbit_r51_c160 bl_160 br_160 wl_51 vdd gnd cell_6t
Xbit_r52_c160 bl_160 br_160 wl_52 vdd gnd cell_6t
Xbit_r53_c160 bl_160 br_160 wl_53 vdd gnd cell_6t
Xbit_r54_c160 bl_160 br_160 wl_54 vdd gnd cell_6t
Xbit_r55_c160 bl_160 br_160 wl_55 vdd gnd cell_6t
Xbit_r56_c160 bl_160 br_160 wl_56 vdd gnd cell_6t
Xbit_r57_c160 bl_160 br_160 wl_57 vdd gnd cell_6t
Xbit_r58_c160 bl_160 br_160 wl_58 vdd gnd cell_6t
Xbit_r59_c160 bl_160 br_160 wl_59 vdd gnd cell_6t
Xbit_r60_c160 bl_160 br_160 wl_60 vdd gnd cell_6t
Xbit_r61_c160 bl_160 br_160 wl_61 vdd gnd cell_6t
Xbit_r62_c160 bl_160 br_160 wl_62 vdd gnd cell_6t
Xbit_r63_c160 bl_160 br_160 wl_63 vdd gnd cell_6t
Xbit_r64_c160 bl_160 br_160 wl_64 vdd gnd cell_6t
Xbit_r65_c160 bl_160 br_160 wl_65 vdd gnd cell_6t
Xbit_r66_c160 bl_160 br_160 wl_66 vdd gnd cell_6t
Xbit_r67_c160 bl_160 br_160 wl_67 vdd gnd cell_6t
Xbit_r68_c160 bl_160 br_160 wl_68 vdd gnd cell_6t
Xbit_r69_c160 bl_160 br_160 wl_69 vdd gnd cell_6t
Xbit_r70_c160 bl_160 br_160 wl_70 vdd gnd cell_6t
Xbit_r71_c160 bl_160 br_160 wl_71 vdd gnd cell_6t
Xbit_r72_c160 bl_160 br_160 wl_72 vdd gnd cell_6t
Xbit_r73_c160 bl_160 br_160 wl_73 vdd gnd cell_6t
Xbit_r74_c160 bl_160 br_160 wl_74 vdd gnd cell_6t
Xbit_r75_c160 bl_160 br_160 wl_75 vdd gnd cell_6t
Xbit_r76_c160 bl_160 br_160 wl_76 vdd gnd cell_6t
Xbit_r77_c160 bl_160 br_160 wl_77 vdd gnd cell_6t
Xbit_r78_c160 bl_160 br_160 wl_78 vdd gnd cell_6t
Xbit_r79_c160 bl_160 br_160 wl_79 vdd gnd cell_6t
Xbit_r80_c160 bl_160 br_160 wl_80 vdd gnd cell_6t
Xbit_r81_c160 bl_160 br_160 wl_81 vdd gnd cell_6t
Xbit_r82_c160 bl_160 br_160 wl_82 vdd gnd cell_6t
Xbit_r83_c160 bl_160 br_160 wl_83 vdd gnd cell_6t
Xbit_r84_c160 bl_160 br_160 wl_84 vdd gnd cell_6t
Xbit_r85_c160 bl_160 br_160 wl_85 vdd gnd cell_6t
Xbit_r86_c160 bl_160 br_160 wl_86 vdd gnd cell_6t
Xbit_r87_c160 bl_160 br_160 wl_87 vdd gnd cell_6t
Xbit_r88_c160 bl_160 br_160 wl_88 vdd gnd cell_6t
Xbit_r89_c160 bl_160 br_160 wl_89 vdd gnd cell_6t
Xbit_r90_c160 bl_160 br_160 wl_90 vdd gnd cell_6t
Xbit_r91_c160 bl_160 br_160 wl_91 vdd gnd cell_6t
Xbit_r92_c160 bl_160 br_160 wl_92 vdd gnd cell_6t
Xbit_r93_c160 bl_160 br_160 wl_93 vdd gnd cell_6t
Xbit_r94_c160 bl_160 br_160 wl_94 vdd gnd cell_6t
Xbit_r95_c160 bl_160 br_160 wl_95 vdd gnd cell_6t
Xbit_r96_c160 bl_160 br_160 wl_96 vdd gnd cell_6t
Xbit_r97_c160 bl_160 br_160 wl_97 vdd gnd cell_6t
Xbit_r98_c160 bl_160 br_160 wl_98 vdd gnd cell_6t
Xbit_r99_c160 bl_160 br_160 wl_99 vdd gnd cell_6t
Xbit_r100_c160 bl_160 br_160 wl_100 vdd gnd cell_6t
Xbit_r101_c160 bl_160 br_160 wl_101 vdd gnd cell_6t
Xbit_r102_c160 bl_160 br_160 wl_102 vdd gnd cell_6t
Xbit_r103_c160 bl_160 br_160 wl_103 vdd gnd cell_6t
Xbit_r104_c160 bl_160 br_160 wl_104 vdd gnd cell_6t
Xbit_r105_c160 bl_160 br_160 wl_105 vdd gnd cell_6t
Xbit_r106_c160 bl_160 br_160 wl_106 vdd gnd cell_6t
Xbit_r107_c160 bl_160 br_160 wl_107 vdd gnd cell_6t
Xbit_r108_c160 bl_160 br_160 wl_108 vdd gnd cell_6t
Xbit_r109_c160 bl_160 br_160 wl_109 vdd gnd cell_6t
Xbit_r110_c160 bl_160 br_160 wl_110 vdd gnd cell_6t
Xbit_r111_c160 bl_160 br_160 wl_111 vdd gnd cell_6t
Xbit_r112_c160 bl_160 br_160 wl_112 vdd gnd cell_6t
Xbit_r113_c160 bl_160 br_160 wl_113 vdd gnd cell_6t
Xbit_r114_c160 bl_160 br_160 wl_114 vdd gnd cell_6t
Xbit_r115_c160 bl_160 br_160 wl_115 vdd gnd cell_6t
Xbit_r116_c160 bl_160 br_160 wl_116 vdd gnd cell_6t
Xbit_r117_c160 bl_160 br_160 wl_117 vdd gnd cell_6t
Xbit_r118_c160 bl_160 br_160 wl_118 vdd gnd cell_6t
Xbit_r119_c160 bl_160 br_160 wl_119 vdd gnd cell_6t
Xbit_r120_c160 bl_160 br_160 wl_120 vdd gnd cell_6t
Xbit_r121_c160 bl_160 br_160 wl_121 vdd gnd cell_6t
Xbit_r122_c160 bl_160 br_160 wl_122 vdd gnd cell_6t
Xbit_r123_c160 bl_160 br_160 wl_123 vdd gnd cell_6t
Xbit_r124_c160 bl_160 br_160 wl_124 vdd gnd cell_6t
Xbit_r125_c160 bl_160 br_160 wl_125 vdd gnd cell_6t
Xbit_r126_c160 bl_160 br_160 wl_126 vdd gnd cell_6t
Xbit_r127_c160 bl_160 br_160 wl_127 vdd gnd cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd cell_6t
Xbit_r1_c161 bl_161 br_161 wl_1 vdd gnd cell_6t
Xbit_r2_c161 bl_161 br_161 wl_2 vdd gnd cell_6t
Xbit_r3_c161 bl_161 br_161 wl_3 vdd gnd cell_6t
Xbit_r4_c161 bl_161 br_161 wl_4 vdd gnd cell_6t
Xbit_r5_c161 bl_161 br_161 wl_5 vdd gnd cell_6t
Xbit_r6_c161 bl_161 br_161 wl_6 vdd gnd cell_6t
Xbit_r7_c161 bl_161 br_161 wl_7 vdd gnd cell_6t
Xbit_r8_c161 bl_161 br_161 wl_8 vdd gnd cell_6t
Xbit_r9_c161 bl_161 br_161 wl_9 vdd gnd cell_6t
Xbit_r10_c161 bl_161 br_161 wl_10 vdd gnd cell_6t
Xbit_r11_c161 bl_161 br_161 wl_11 vdd gnd cell_6t
Xbit_r12_c161 bl_161 br_161 wl_12 vdd gnd cell_6t
Xbit_r13_c161 bl_161 br_161 wl_13 vdd gnd cell_6t
Xbit_r14_c161 bl_161 br_161 wl_14 vdd gnd cell_6t
Xbit_r15_c161 bl_161 br_161 wl_15 vdd gnd cell_6t
Xbit_r16_c161 bl_161 br_161 wl_16 vdd gnd cell_6t
Xbit_r17_c161 bl_161 br_161 wl_17 vdd gnd cell_6t
Xbit_r18_c161 bl_161 br_161 wl_18 vdd gnd cell_6t
Xbit_r19_c161 bl_161 br_161 wl_19 vdd gnd cell_6t
Xbit_r20_c161 bl_161 br_161 wl_20 vdd gnd cell_6t
Xbit_r21_c161 bl_161 br_161 wl_21 vdd gnd cell_6t
Xbit_r22_c161 bl_161 br_161 wl_22 vdd gnd cell_6t
Xbit_r23_c161 bl_161 br_161 wl_23 vdd gnd cell_6t
Xbit_r24_c161 bl_161 br_161 wl_24 vdd gnd cell_6t
Xbit_r25_c161 bl_161 br_161 wl_25 vdd gnd cell_6t
Xbit_r26_c161 bl_161 br_161 wl_26 vdd gnd cell_6t
Xbit_r27_c161 bl_161 br_161 wl_27 vdd gnd cell_6t
Xbit_r28_c161 bl_161 br_161 wl_28 vdd gnd cell_6t
Xbit_r29_c161 bl_161 br_161 wl_29 vdd gnd cell_6t
Xbit_r30_c161 bl_161 br_161 wl_30 vdd gnd cell_6t
Xbit_r31_c161 bl_161 br_161 wl_31 vdd gnd cell_6t
Xbit_r32_c161 bl_161 br_161 wl_32 vdd gnd cell_6t
Xbit_r33_c161 bl_161 br_161 wl_33 vdd gnd cell_6t
Xbit_r34_c161 bl_161 br_161 wl_34 vdd gnd cell_6t
Xbit_r35_c161 bl_161 br_161 wl_35 vdd gnd cell_6t
Xbit_r36_c161 bl_161 br_161 wl_36 vdd gnd cell_6t
Xbit_r37_c161 bl_161 br_161 wl_37 vdd gnd cell_6t
Xbit_r38_c161 bl_161 br_161 wl_38 vdd gnd cell_6t
Xbit_r39_c161 bl_161 br_161 wl_39 vdd gnd cell_6t
Xbit_r40_c161 bl_161 br_161 wl_40 vdd gnd cell_6t
Xbit_r41_c161 bl_161 br_161 wl_41 vdd gnd cell_6t
Xbit_r42_c161 bl_161 br_161 wl_42 vdd gnd cell_6t
Xbit_r43_c161 bl_161 br_161 wl_43 vdd gnd cell_6t
Xbit_r44_c161 bl_161 br_161 wl_44 vdd gnd cell_6t
Xbit_r45_c161 bl_161 br_161 wl_45 vdd gnd cell_6t
Xbit_r46_c161 bl_161 br_161 wl_46 vdd gnd cell_6t
Xbit_r47_c161 bl_161 br_161 wl_47 vdd gnd cell_6t
Xbit_r48_c161 bl_161 br_161 wl_48 vdd gnd cell_6t
Xbit_r49_c161 bl_161 br_161 wl_49 vdd gnd cell_6t
Xbit_r50_c161 bl_161 br_161 wl_50 vdd gnd cell_6t
Xbit_r51_c161 bl_161 br_161 wl_51 vdd gnd cell_6t
Xbit_r52_c161 bl_161 br_161 wl_52 vdd gnd cell_6t
Xbit_r53_c161 bl_161 br_161 wl_53 vdd gnd cell_6t
Xbit_r54_c161 bl_161 br_161 wl_54 vdd gnd cell_6t
Xbit_r55_c161 bl_161 br_161 wl_55 vdd gnd cell_6t
Xbit_r56_c161 bl_161 br_161 wl_56 vdd gnd cell_6t
Xbit_r57_c161 bl_161 br_161 wl_57 vdd gnd cell_6t
Xbit_r58_c161 bl_161 br_161 wl_58 vdd gnd cell_6t
Xbit_r59_c161 bl_161 br_161 wl_59 vdd gnd cell_6t
Xbit_r60_c161 bl_161 br_161 wl_60 vdd gnd cell_6t
Xbit_r61_c161 bl_161 br_161 wl_61 vdd gnd cell_6t
Xbit_r62_c161 bl_161 br_161 wl_62 vdd gnd cell_6t
Xbit_r63_c161 bl_161 br_161 wl_63 vdd gnd cell_6t
Xbit_r64_c161 bl_161 br_161 wl_64 vdd gnd cell_6t
Xbit_r65_c161 bl_161 br_161 wl_65 vdd gnd cell_6t
Xbit_r66_c161 bl_161 br_161 wl_66 vdd gnd cell_6t
Xbit_r67_c161 bl_161 br_161 wl_67 vdd gnd cell_6t
Xbit_r68_c161 bl_161 br_161 wl_68 vdd gnd cell_6t
Xbit_r69_c161 bl_161 br_161 wl_69 vdd gnd cell_6t
Xbit_r70_c161 bl_161 br_161 wl_70 vdd gnd cell_6t
Xbit_r71_c161 bl_161 br_161 wl_71 vdd gnd cell_6t
Xbit_r72_c161 bl_161 br_161 wl_72 vdd gnd cell_6t
Xbit_r73_c161 bl_161 br_161 wl_73 vdd gnd cell_6t
Xbit_r74_c161 bl_161 br_161 wl_74 vdd gnd cell_6t
Xbit_r75_c161 bl_161 br_161 wl_75 vdd gnd cell_6t
Xbit_r76_c161 bl_161 br_161 wl_76 vdd gnd cell_6t
Xbit_r77_c161 bl_161 br_161 wl_77 vdd gnd cell_6t
Xbit_r78_c161 bl_161 br_161 wl_78 vdd gnd cell_6t
Xbit_r79_c161 bl_161 br_161 wl_79 vdd gnd cell_6t
Xbit_r80_c161 bl_161 br_161 wl_80 vdd gnd cell_6t
Xbit_r81_c161 bl_161 br_161 wl_81 vdd gnd cell_6t
Xbit_r82_c161 bl_161 br_161 wl_82 vdd gnd cell_6t
Xbit_r83_c161 bl_161 br_161 wl_83 vdd gnd cell_6t
Xbit_r84_c161 bl_161 br_161 wl_84 vdd gnd cell_6t
Xbit_r85_c161 bl_161 br_161 wl_85 vdd gnd cell_6t
Xbit_r86_c161 bl_161 br_161 wl_86 vdd gnd cell_6t
Xbit_r87_c161 bl_161 br_161 wl_87 vdd gnd cell_6t
Xbit_r88_c161 bl_161 br_161 wl_88 vdd gnd cell_6t
Xbit_r89_c161 bl_161 br_161 wl_89 vdd gnd cell_6t
Xbit_r90_c161 bl_161 br_161 wl_90 vdd gnd cell_6t
Xbit_r91_c161 bl_161 br_161 wl_91 vdd gnd cell_6t
Xbit_r92_c161 bl_161 br_161 wl_92 vdd gnd cell_6t
Xbit_r93_c161 bl_161 br_161 wl_93 vdd gnd cell_6t
Xbit_r94_c161 bl_161 br_161 wl_94 vdd gnd cell_6t
Xbit_r95_c161 bl_161 br_161 wl_95 vdd gnd cell_6t
Xbit_r96_c161 bl_161 br_161 wl_96 vdd gnd cell_6t
Xbit_r97_c161 bl_161 br_161 wl_97 vdd gnd cell_6t
Xbit_r98_c161 bl_161 br_161 wl_98 vdd gnd cell_6t
Xbit_r99_c161 bl_161 br_161 wl_99 vdd gnd cell_6t
Xbit_r100_c161 bl_161 br_161 wl_100 vdd gnd cell_6t
Xbit_r101_c161 bl_161 br_161 wl_101 vdd gnd cell_6t
Xbit_r102_c161 bl_161 br_161 wl_102 vdd gnd cell_6t
Xbit_r103_c161 bl_161 br_161 wl_103 vdd gnd cell_6t
Xbit_r104_c161 bl_161 br_161 wl_104 vdd gnd cell_6t
Xbit_r105_c161 bl_161 br_161 wl_105 vdd gnd cell_6t
Xbit_r106_c161 bl_161 br_161 wl_106 vdd gnd cell_6t
Xbit_r107_c161 bl_161 br_161 wl_107 vdd gnd cell_6t
Xbit_r108_c161 bl_161 br_161 wl_108 vdd gnd cell_6t
Xbit_r109_c161 bl_161 br_161 wl_109 vdd gnd cell_6t
Xbit_r110_c161 bl_161 br_161 wl_110 vdd gnd cell_6t
Xbit_r111_c161 bl_161 br_161 wl_111 vdd gnd cell_6t
Xbit_r112_c161 bl_161 br_161 wl_112 vdd gnd cell_6t
Xbit_r113_c161 bl_161 br_161 wl_113 vdd gnd cell_6t
Xbit_r114_c161 bl_161 br_161 wl_114 vdd gnd cell_6t
Xbit_r115_c161 bl_161 br_161 wl_115 vdd gnd cell_6t
Xbit_r116_c161 bl_161 br_161 wl_116 vdd gnd cell_6t
Xbit_r117_c161 bl_161 br_161 wl_117 vdd gnd cell_6t
Xbit_r118_c161 bl_161 br_161 wl_118 vdd gnd cell_6t
Xbit_r119_c161 bl_161 br_161 wl_119 vdd gnd cell_6t
Xbit_r120_c161 bl_161 br_161 wl_120 vdd gnd cell_6t
Xbit_r121_c161 bl_161 br_161 wl_121 vdd gnd cell_6t
Xbit_r122_c161 bl_161 br_161 wl_122 vdd gnd cell_6t
Xbit_r123_c161 bl_161 br_161 wl_123 vdd gnd cell_6t
Xbit_r124_c161 bl_161 br_161 wl_124 vdd gnd cell_6t
Xbit_r125_c161 bl_161 br_161 wl_125 vdd gnd cell_6t
Xbit_r126_c161 bl_161 br_161 wl_126 vdd gnd cell_6t
Xbit_r127_c161 bl_161 br_161 wl_127 vdd gnd cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd cell_6t
Xbit_r1_c162 bl_162 br_162 wl_1 vdd gnd cell_6t
Xbit_r2_c162 bl_162 br_162 wl_2 vdd gnd cell_6t
Xbit_r3_c162 bl_162 br_162 wl_3 vdd gnd cell_6t
Xbit_r4_c162 bl_162 br_162 wl_4 vdd gnd cell_6t
Xbit_r5_c162 bl_162 br_162 wl_5 vdd gnd cell_6t
Xbit_r6_c162 bl_162 br_162 wl_6 vdd gnd cell_6t
Xbit_r7_c162 bl_162 br_162 wl_7 vdd gnd cell_6t
Xbit_r8_c162 bl_162 br_162 wl_8 vdd gnd cell_6t
Xbit_r9_c162 bl_162 br_162 wl_9 vdd gnd cell_6t
Xbit_r10_c162 bl_162 br_162 wl_10 vdd gnd cell_6t
Xbit_r11_c162 bl_162 br_162 wl_11 vdd gnd cell_6t
Xbit_r12_c162 bl_162 br_162 wl_12 vdd gnd cell_6t
Xbit_r13_c162 bl_162 br_162 wl_13 vdd gnd cell_6t
Xbit_r14_c162 bl_162 br_162 wl_14 vdd gnd cell_6t
Xbit_r15_c162 bl_162 br_162 wl_15 vdd gnd cell_6t
Xbit_r16_c162 bl_162 br_162 wl_16 vdd gnd cell_6t
Xbit_r17_c162 bl_162 br_162 wl_17 vdd gnd cell_6t
Xbit_r18_c162 bl_162 br_162 wl_18 vdd gnd cell_6t
Xbit_r19_c162 bl_162 br_162 wl_19 vdd gnd cell_6t
Xbit_r20_c162 bl_162 br_162 wl_20 vdd gnd cell_6t
Xbit_r21_c162 bl_162 br_162 wl_21 vdd gnd cell_6t
Xbit_r22_c162 bl_162 br_162 wl_22 vdd gnd cell_6t
Xbit_r23_c162 bl_162 br_162 wl_23 vdd gnd cell_6t
Xbit_r24_c162 bl_162 br_162 wl_24 vdd gnd cell_6t
Xbit_r25_c162 bl_162 br_162 wl_25 vdd gnd cell_6t
Xbit_r26_c162 bl_162 br_162 wl_26 vdd gnd cell_6t
Xbit_r27_c162 bl_162 br_162 wl_27 vdd gnd cell_6t
Xbit_r28_c162 bl_162 br_162 wl_28 vdd gnd cell_6t
Xbit_r29_c162 bl_162 br_162 wl_29 vdd gnd cell_6t
Xbit_r30_c162 bl_162 br_162 wl_30 vdd gnd cell_6t
Xbit_r31_c162 bl_162 br_162 wl_31 vdd gnd cell_6t
Xbit_r32_c162 bl_162 br_162 wl_32 vdd gnd cell_6t
Xbit_r33_c162 bl_162 br_162 wl_33 vdd gnd cell_6t
Xbit_r34_c162 bl_162 br_162 wl_34 vdd gnd cell_6t
Xbit_r35_c162 bl_162 br_162 wl_35 vdd gnd cell_6t
Xbit_r36_c162 bl_162 br_162 wl_36 vdd gnd cell_6t
Xbit_r37_c162 bl_162 br_162 wl_37 vdd gnd cell_6t
Xbit_r38_c162 bl_162 br_162 wl_38 vdd gnd cell_6t
Xbit_r39_c162 bl_162 br_162 wl_39 vdd gnd cell_6t
Xbit_r40_c162 bl_162 br_162 wl_40 vdd gnd cell_6t
Xbit_r41_c162 bl_162 br_162 wl_41 vdd gnd cell_6t
Xbit_r42_c162 bl_162 br_162 wl_42 vdd gnd cell_6t
Xbit_r43_c162 bl_162 br_162 wl_43 vdd gnd cell_6t
Xbit_r44_c162 bl_162 br_162 wl_44 vdd gnd cell_6t
Xbit_r45_c162 bl_162 br_162 wl_45 vdd gnd cell_6t
Xbit_r46_c162 bl_162 br_162 wl_46 vdd gnd cell_6t
Xbit_r47_c162 bl_162 br_162 wl_47 vdd gnd cell_6t
Xbit_r48_c162 bl_162 br_162 wl_48 vdd gnd cell_6t
Xbit_r49_c162 bl_162 br_162 wl_49 vdd gnd cell_6t
Xbit_r50_c162 bl_162 br_162 wl_50 vdd gnd cell_6t
Xbit_r51_c162 bl_162 br_162 wl_51 vdd gnd cell_6t
Xbit_r52_c162 bl_162 br_162 wl_52 vdd gnd cell_6t
Xbit_r53_c162 bl_162 br_162 wl_53 vdd gnd cell_6t
Xbit_r54_c162 bl_162 br_162 wl_54 vdd gnd cell_6t
Xbit_r55_c162 bl_162 br_162 wl_55 vdd gnd cell_6t
Xbit_r56_c162 bl_162 br_162 wl_56 vdd gnd cell_6t
Xbit_r57_c162 bl_162 br_162 wl_57 vdd gnd cell_6t
Xbit_r58_c162 bl_162 br_162 wl_58 vdd gnd cell_6t
Xbit_r59_c162 bl_162 br_162 wl_59 vdd gnd cell_6t
Xbit_r60_c162 bl_162 br_162 wl_60 vdd gnd cell_6t
Xbit_r61_c162 bl_162 br_162 wl_61 vdd gnd cell_6t
Xbit_r62_c162 bl_162 br_162 wl_62 vdd gnd cell_6t
Xbit_r63_c162 bl_162 br_162 wl_63 vdd gnd cell_6t
Xbit_r64_c162 bl_162 br_162 wl_64 vdd gnd cell_6t
Xbit_r65_c162 bl_162 br_162 wl_65 vdd gnd cell_6t
Xbit_r66_c162 bl_162 br_162 wl_66 vdd gnd cell_6t
Xbit_r67_c162 bl_162 br_162 wl_67 vdd gnd cell_6t
Xbit_r68_c162 bl_162 br_162 wl_68 vdd gnd cell_6t
Xbit_r69_c162 bl_162 br_162 wl_69 vdd gnd cell_6t
Xbit_r70_c162 bl_162 br_162 wl_70 vdd gnd cell_6t
Xbit_r71_c162 bl_162 br_162 wl_71 vdd gnd cell_6t
Xbit_r72_c162 bl_162 br_162 wl_72 vdd gnd cell_6t
Xbit_r73_c162 bl_162 br_162 wl_73 vdd gnd cell_6t
Xbit_r74_c162 bl_162 br_162 wl_74 vdd gnd cell_6t
Xbit_r75_c162 bl_162 br_162 wl_75 vdd gnd cell_6t
Xbit_r76_c162 bl_162 br_162 wl_76 vdd gnd cell_6t
Xbit_r77_c162 bl_162 br_162 wl_77 vdd gnd cell_6t
Xbit_r78_c162 bl_162 br_162 wl_78 vdd gnd cell_6t
Xbit_r79_c162 bl_162 br_162 wl_79 vdd gnd cell_6t
Xbit_r80_c162 bl_162 br_162 wl_80 vdd gnd cell_6t
Xbit_r81_c162 bl_162 br_162 wl_81 vdd gnd cell_6t
Xbit_r82_c162 bl_162 br_162 wl_82 vdd gnd cell_6t
Xbit_r83_c162 bl_162 br_162 wl_83 vdd gnd cell_6t
Xbit_r84_c162 bl_162 br_162 wl_84 vdd gnd cell_6t
Xbit_r85_c162 bl_162 br_162 wl_85 vdd gnd cell_6t
Xbit_r86_c162 bl_162 br_162 wl_86 vdd gnd cell_6t
Xbit_r87_c162 bl_162 br_162 wl_87 vdd gnd cell_6t
Xbit_r88_c162 bl_162 br_162 wl_88 vdd gnd cell_6t
Xbit_r89_c162 bl_162 br_162 wl_89 vdd gnd cell_6t
Xbit_r90_c162 bl_162 br_162 wl_90 vdd gnd cell_6t
Xbit_r91_c162 bl_162 br_162 wl_91 vdd gnd cell_6t
Xbit_r92_c162 bl_162 br_162 wl_92 vdd gnd cell_6t
Xbit_r93_c162 bl_162 br_162 wl_93 vdd gnd cell_6t
Xbit_r94_c162 bl_162 br_162 wl_94 vdd gnd cell_6t
Xbit_r95_c162 bl_162 br_162 wl_95 vdd gnd cell_6t
Xbit_r96_c162 bl_162 br_162 wl_96 vdd gnd cell_6t
Xbit_r97_c162 bl_162 br_162 wl_97 vdd gnd cell_6t
Xbit_r98_c162 bl_162 br_162 wl_98 vdd gnd cell_6t
Xbit_r99_c162 bl_162 br_162 wl_99 vdd gnd cell_6t
Xbit_r100_c162 bl_162 br_162 wl_100 vdd gnd cell_6t
Xbit_r101_c162 bl_162 br_162 wl_101 vdd gnd cell_6t
Xbit_r102_c162 bl_162 br_162 wl_102 vdd gnd cell_6t
Xbit_r103_c162 bl_162 br_162 wl_103 vdd gnd cell_6t
Xbit_r104_c162 bl_162 br_162 wl_104 vdd gnd cell_6t
Xbit_r105_c162 bl_162 br_162 wl_105 vdd gnd cell_6t
Xbit_r106_c162 bl_162 br_162 wl_106 vdd gnd cell_6t
Xbit_r107_c162 bl_162 br_162 wl_107 vdd gnd cell_6t
Xbit_r108_c162 bl_162 br_162 wl_108 vdd gnd cell_6t
Xbit_r109_c162 bl_162 br_162 wl_109 vdd gnd cell_6t
Xbit_r110_c162 bl_162 br_162 wl_110 vdd gnd cell_6t
Xbit_r111_c162 bl_162 br_162 wl_111 vdd gnd cell_6t
Xbit_r112_c162 bl_162 br_162 wl_112 vdd gnd cell_6t
Xbit_r113_c162 bl_162 br_162 wl_113 vdd gnd cell_6t
Xbit_r114_c162 bl_162 br_162 wl_114 vdd gnd cell_6t
Xbit_r115_c162 bl_162 br_162 wl_115 vdd gnd cell_6t
Xbit_r116_c162 bl_162 br_162 wl_116 vdd gnd cell_6t
Xbit_r117_c162 bl_162 br_162 wl_117 vdd gnd cell_6t
Xbit_r118_c162 bl_162 br_162 wl_118 vdd gnd cell_6t
Xbit_r119_c162 bl_162 br_162 wl_119 vdd gnd cell_6t
Xbit_r120_c162 bl_162 br_162 wl_120 vdd gnd cell_6t
Xbit_r121_c162 bl_162 br_162 wl_121 vdd gnd cell_6t
Xbit_r122_c162 bl_162 br_162 wl_122 vdd gnd cell_6t
Xbit_r123_c162 bl_162 br_162 wl_123 vdd gnd cell_6t
Xbit_r124_c162 bl_162 br_162 wl_124 vdd gnd cell_6t
Xbit_r125_c162 bl_162 br_162 wl_125 vdd gnd cell_6t
Xbit_r126_c162 bl_162 br_162 wl_126 vdd gnd cell_6t
Xbit_r127_c162 bl_162 br_162 wl_127 vdd gnd cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd cell_6t
Xbit_r1_c163 bl_163 br_163 wl_1 vdd gnd cell_6t
Xbit_r2_c163 bl_163 br_163 wl_2 vdd gnd cell_6t
Xbit_r3_c163 bl_163 br_163 wl_3 vdd gnd cell_6t
Xbit_r4_c163 bl_163 br_163 wl_4 vdd gnd cell_6t
Xbit_r5_c163 bl_163 br_163 wl_5 vdd gnd cell_6t
Xbit_r6_c163 bl_163 br_163 wl_6 vdd gnd cell_6t
Xbit_r7_c163 bl_163 br_163 wl_7 vdd gnd cell_6t
Xbit_r8_c163 bl_163 br_163 wl_8 vdd gnd cell_6t
Xbit_r9_c163 bl_163 br_163 wl_9 vdd gnd cell_6t
Xbit_r10_c163 bl_163 br_163 wl_10 vdd gnd cell_6t
Xbit_r11_c163 bl_163 br_163 wl_11 vdd gnd cell_6t
Xbit_r12_c163 bl_163 br_163 wl_12 vdd gnd cell_6t
Xbit_r13_c163 bl_163 br_163 wl_13 vdd gnd cell_6t
Xbit_r14_c163 bl_163 br_163 wl_14 vdd gnd cell_6t
Xbit_r15_c163 bl_163 br_163 wl_15 vdd gnd cell_6t
Xbit_r16_c163 bl_163 br_163 wl_16 vdd gnd cell_6t
Xbit_r17_c163 bl_163 br_163 wl_17 vdd gnd cell_6t
Xbit_r18_c163 bl_163 br_163 wl_18 vdd gnd cell_6t
Xbit_r19_c163 bl_163 br_163 wl_19 vdd gnd cell_6t
Xbit_r20_c163 bl_163 br_163 wl_20 vdd gnd cell_6t
Xbit_r21_c163 bl_163 br_163 wl_21 vdd gnd cell_6t
Xbit_r22_c163 bl_163 br_163 wl_22 vdd gnd cell_6t
Xbit_r23_c163 bl_163 br_163 wl_23 vdd gnd cell_6t
Xbit_r24_c163 bl_163 br_163 wl_24 vdd gnd cell_6t
Xbit_r25_c163 bl_163 br_163 wl_25 vdd gnd cell_6t
Xbit_r26_c163 bl_163 br_163 wl_26 vdd gnd cell_6t
Xbit_r27_c163 bl_163 br_163 wl_27 vdd gnd cell_6t
Xbit_r28_c163 bl_163 br_163 wl_28 vdd gnd cell_6t
Xbit_r29_c163 bl_163 br_163 wl_29 vdd gnd cell_6t
Xbit_r30_c163 bl_163 br_163 wl_30 vdd gnd cell_6t
Xbit_r31_c163 bl_163 br_163 wl_31 vdd gnd cell_6t
Xbit_r32_c163 bl_163 br_163 wl_32 vdd gnd cell_6t
Xbit_r33_c163 bl_163 br_163 wl_33 vdd gnd cell_6t
Xbit_r34_c163 bl_163 br_163 wl_34 vdd gnd cell_6t
Xbit_r35_c163 bl_163 br_163 wl_35 vdd gnd cell_6t
Xbit_r36_c163 bl_163 br_163 wl_36 vdd gnd cell_6t
Xbit_r37_c163 bl_163 br_163 wl_37 vdd gnd cell_6t
Xbit_r38_c163 bl_163 br_163 wl_38 vdd gnd cell_6t
Xbit_r39_c163 bl_163 br_163 wl_39 vdd gnd cell_6t
Xbit_r40_c163 bl_163 br_163 wl_40 vdd gnd cell_6t
Xbit_r41_c163 bl_163 br_163 wl_41 vdd gnd cell_6t
Xbit_r42_c163 bl_163 br_163 wl_42 vdd gnd cell_6t
Xbit_r43_c163 bl_163 br_163 wl_43 vdd gnd cell_6t
Xbit_r44_c163 bl_163 br_163 wl_44 vdd gnd cell_6t
Xbit_r45_c163 bl_163 br_163 wl_45 vdd gnd cell_6t
Xbit_r46_c163 bl_163 br_163 wl_46 vdd gnd cell_6t
Xbit_r47_c163 bl_163 br_163 wl_47 vdd gnd cell_6t
Xbit_r48_c163 bl_163 br_163 wl_48 vdd gnd cell_6t
Xbit_r49_c163 bl_163 br_163 wl_49 vdd gnd cell_6t
Xbit_r50_c163 bl_163 br_163 wl_50 vdd gnd cell_6t
Xbit_r51_c163 bl_163 br_163 wl_51 vdd gnd cell_6t
Xbit_r52_c163 bl_163 br_163 wl_52 vdd gnd cell_6t
Xbit_r53_c163 bl_163 br_163 wl_53 vdd gnd cell_6t
Xbit_r54_c163 bl_163 br_163 wl_54 vdd gnd cell_6t
Xbit_r55_c163 bl_163 br_163 wl_55 vdd gnd cell_6t
Xbit_r56_c163 bl_163 br_163 wl_56 vdd gnd cell_6t
Xbit_r57_c163 bl_163 br_163 wl_57 vdd gnd cell_6t
Xbit_r58_c163 bl_163 br_163 wl_58 vdd gnd cell_6t
Xbit_r59_c163 bl_163 br_163 wl_59 vdd gnd cell_6t
Xbit_r60_c163 bl_163 br_163 wl_60 vdd gnd cell_6t
Xbit_r61_c163 bl_163 br_163 wl_61 vdd gnd cell_6t
Xbit_r62_c163 bl_163 br_163 wl_62 vdd gnd cell_6t
Xbit_r63_c163 bl_163 br_163 wl_63 vdd gnd cell_6t
Xbit_r64_c163 bl_163 br_163 wl_64 vdd gnd cell_6t
Xbit_r65_c163 bl_163 br_163 wl_65 vdd gnd cell_6t
Xbit_r66_c163 bl_163 br_163 wl_66 vdd gnd cell_6t
Xbit_r67_c163 bl_163 br_163 wl_67 vdd gnd cell_6t
Xbit_r68_c163 bl_163 br_163 wl_68 vdd gnd cell_6t
Xbit_r69_c163 bl_163 br_163 wl_69 vdd gnd cell_6t
Xbit_r70_c163 bl_163 br_163 wl_70 vdd gnd cell_6t
Xbit_r71_c163 bl_163 br_163 wl_71 vdd gnd cell_6t
Xbit_r72_c163 bl_163 br_163 wl_72 vdd gnd cell_6t
Xbit_r73_c163 bl_163 br_163 wl_73 vdd gnd cell_6t
Xbit_r74_c163 bl_163 br_163 wl_74 vdd gnd cell_6t
Xbit_r75_c163 bl_163 br_163 wl_75 vdd gnd cell_6t
Xbit_r76_c163 bl_163 br_163 wl_76 vdd gnd cell_6t
Xbit_r77_c163 bl_163 br_163 wl_77 vdd gnd cell_6t
Xbit_r78_c163 bl_163 br_163 wl_78 vdd gnd cell_6t
Xbit_r79_c163 bl_163 br_163 wl_79 vdd gnd cell_6t
Xbit_r80_c163 bl_163 br_163 wl_80 vdd gnd cell_6t
Xbit_r81_c163 bl_163 br_163 wl_81 vdd gnd cell_6t
Xbit_r82_c163 bl_163 br_163 wl_82 vdd gnd cell_6t
Xbit_r83_c163 bl_163 br_163 wl_83 vdd gnd cell_6t
Xbit_r84_c163 bl_163 br_163 wl_84 vdd gnd cell_6t
Xbit_r85_c163 bl_163 br_163 wl_85 vdd gnd cell_6t
Xbit_r86_c163 bl_163 br_163 wl_86 vdd gnd cell_6t
Xbit_r87_c163 bl_163 br_163 wl_87 vdd gnd cell_6t
Xbit_r88_c163 bl_163 br_163 wl_88 vdd gnd cell_6t
Xbit_r89_c163 bl_163 br_163 wl_89 vdd gnd cell_6t
Xbit_r90_c163 bl_163 br_163 wl_90 vdd gnd cell_6t
Xbit_r91_c163 bl_163 br_163 wl_91 vdd gnd cell_6t
Xbit_r92_c163 bl_163 br_163 wl_92 vdd gnd cell_6t
Xbit_r93_c163 bl_163 br_163 wl_93 vdd gnd cell_6t
Xbit_r94_c163 bl_163 br_163 wl_94 vdd gnd cell_6t
Xbit_r95_c163 bl_163 br_163 wl_95 vdd gnd cell_6t
Xbit_r96_c163 bl_163 br_163 wl_96 vdd gnd cell_6t
Xbit_r97_c163 bl_163 br_163 wl_97 vdd gnd cell_6t
Xbit_r98_c163 bl_163 br_163 wl_98 vdd gnd cell_6t
Xbit_r99_c163 bl_163 br_163 wl_99 vdd gnd cell_6t
Xbit_r100_c163 bl_163 br_163 wl_100 vdd gnd cell_6t
Xbit_r101_c163 bl_163 br_163 wl_101 vdd gnd cell_6t
Xbit_r102_c163 bl_163 br_163 wl_102 vdd gnd cell_6t
Xbit_r103_c163 bl_163 br_163 wl_103 vdd gnd cell_6t
Xbit_r104_c163 bl_163 br_163 wl_104 vdd gnd cell_6t
Xbit_r105_c163 bl_163 br_163 wl_105 vdd gnd cell_6t
Xbit_r106_c163 bl_163 br_163 wl_106 vdd gnd cell_6t
Xbit_r107_c163 bl_163 br_163 wl_107 vdd gnd cell_6t
Xbit_r108_c163 bl_163 br_163 wl_108 vdd gnd cell_6t
Xbit_r109_c163 bl_163 br_163 wl_109 vdd gnd cell_6t
Xbit_r110_c163 bl_163 br_163 wl_110 vdd gnd cell_6t
Xbit_r111_c163 bl_163 br_163 wl_111 vdd gnd cell_6t
Xbit_r112_c163 bl_163 br_163 wl_112 vdd gnd cell_6t
Xbit_r113_c163 bl_163 br_163 wl_113 vdd gnd cell_6t
Xbit_r114_c163 bl_163 br_163 wl_114 vdd gnd cell_6t
Xbit_r115_c163 bl_163 br_163 wl_115 vdd gnd cell_6t
Xbit_r116_c163 bl_163 br_163 wl_116 vdd gnd cell_6t
Xbit_r117_c163 bl_163 br_163 wl_117 vdd gnd cell_6t
Xbit_r118_c163 bl_163 br_163 wl_118 vdd gnd cell_6t
Xbit_r119_c163 bl_163 br_163 wl_119 vdd gnd cell_6t
Xbit_r120_c163 bl_163 br_163 wl_120 vdd gnd cell_6t
Xbit_r121_c163 bl_163 br_163 wl_121 vdd gnd cell_6t
Xbit_r122_c163 bl_163 br_163 wl_122 vdd gnd cell_6t
Xbit_r123_c163 bl_163 br_163 wl_123 vdd gnd cell_6t
Xbit_r124_c163 bl_163 br_163 wl_124 vdd gnd cell_6t
Xbit_r125_c163 bl_163 br_163 wl_125 vdd gnd cell_6t
Xbit_r126_c163 bl_163 br_163 wl_126 vdd gnd cell_6t
Xbit_r127_c163 bl_163 br_163 wl_127 vdd gnd cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd cell_6t
Xbit_r1_c164 bl_164 br_164 wl_1 vdd gnd cell_6t
Xbit_r2_c164 bl_164 br_164 wl_2 vdd gnd cell_6t
Xbit_r3_c164 bl_164 br_164 wl_3 vdd gnd cell_6t
Xbit_r4_c164 bl_164 br_164 wl_4 vdd gnd cell_6t
Xbit_r5_c164 bl_164 br_164 wl_5 vdd gnd cell_6t
Xbit_r6_c164 bl_164 br_164 wl_6 vdd gnd cell_6t
Xbit_r7_c164 bl_164 br_164 wl_7 vdd gnd cell_6t
Xbit_r8_c164 bl_164 br_164 wl_8 vdd gnd cell_6t
Xbit_r9_c164 bl_164 br_164 wl_9 vdd gnd cell_6t
Xbit_r10_c164 bl_164 br_164 wl_10 vdd gnd cell_6t
Xbit_r11_c164 bl_164 br_164 wl_11 vdd gnd cell_6t
Xbit_r12_c164 bl_164 br_164 wl_12 vdd gnd cell_6t
Xbit_r13_c164 bl_164 br_164 wl_13 vdd gnd cell_6t
Xbit_r14_c164 bl_164 br_164 wl_14 vdd gnd cell_6t
Xbit_r15_c164 bl_164 br_164 wl_15 vdd gnd cell_6t
Xbit_r16_c164 bl_164 br_164 wl_16 vdd gnd cell_6t
Xbit_r17_c164 bl_164 br_164 wl_17 vdd gnd cell_6t
Xbit_r18_c164 bl_164 br_164 wl_18 vdd gnd cell_6t
Xbit_r19_c164 bl_164 br_164 wl_19 vdd gnd cell_6t
Xbit_r20_c164 bl_164 br_164 wl_20 vdd gnd cell_6t
Xbit_r21_c164 bl_164 br_164 wl_21 vdd gnd cell_6t
Xbit_r22_c164 bl_164 br_164 wl_22 vdd gnd cell_6t
Xbit_r23_c164 bl_164 br_164 wl_23 vdd gnd cell_6t
Xbit_r24_c164 bl_164 br_164 wl_24 vdd gnd cell_6t
Xbit_r25_c164 bl_164 br_164 wl_25 vdd gnd cell_6t
Xbit_r26_c164 bl_164 br_164 wl_26 vdd gnd cell_6t
Xbit_r27_c164 bl_164 br_164 wl_27 vdd gnd cell_6t
Xbit_r28_c164 bl_164 br_164 wl_28 vdd gnd cell_6t
Xbit_r29_c164 bl_164 br_164 wl_29 vdd gnd cell_6t
Xbit_r30_c164 bl_164 br_164 wl_30 vdd gnd cell_6t
Xbit_r31_c164 bl_164 br_164 wl_31 vdd gnd cell_6t
Xbit_r32_c164 bl_164 br_164 wl_32 vdd gnd cell_6t
Xbit_r33_c164 bl_164 br_164 wl_33 vdd gnd cell_6t
Xbit_r34_c164 bl_164 br_164 wl_34 vdd gnd cell_6t
Xbit_r35_c164 bl_164 br_164 wl_35 vdd gnd cell_6t
Xbit_r36_c164 bl_164 br_164 wl_36 vdd gnd cell_6t
Xbit_r37_c164 bl_164 br_164 wl_37 vdd gnd cell_6t
Xbit_r38_c164 bl_164 br_164 wl_38 vdd gnd cell_6t
Xbit_r39_c164 bl_164 br_164 wl_39 vdd gnd cell_6t
Xbit_r40_c164 bl_164 br_164 wl_40 vdd gnd cell_6t
Xbit_r41_c164 bl_164 br_164 wl_41 vdd gnd cell_6t
Xbit_r42_c164 bl_164 br_164 wl_42 vdd gnd cell_6t
Xbit_r43_c164 bl_164 br_164 wl_43 vdd gnd cell_6t
Xbit_r44_c164 bl_164 br_164 wl_44 vdd gnd cell_6t
Xbit_r45_c164 bl_164 br_164 wl_45 vdd gnd cell_6t
Xbit_r46_c164 bl_164 br_164 wl_46 vdd gnd cell_6t
Xbit_r47_c164 bl_164 br_164 wl_47 vdd gnd cell_6t
Xbit_r48_c164 bl_164 br_164 wl_48 vdd gnd cell_6t
Xbit_r49_c164 bl_164 br_164 wl_49 vdd gnd cell_6t
Xbit_r50_c164 bl_164 br_164 wl_50 vdd gnd cell_6t
Xbit_r51_c164 bl_164 br_164 wl_51 vdd gnd cell_6t
Xbit_r52_c164 bl_164 br_164 wl_52 vdd gnd cell_6t
Xbit_r53_c164 bl_164 br_164 wl_53 vdd gnd cell_6t
Xbit_r54_c164 bl_164 br_164 wl_54 vdd gnd cell_6t
Xbit_r55_c164 bl_164 br_164 wl_55 vdd gnd cell_6t
Xbit_r56_c164 bl_164 br_164 wl_56 vdd gnd cell_6t
Xbit_r57_c164 bl_164 br_164 wl_57 vdd gnd cell_6t
Xbit_r58_c164 bl_164 br_164 wl_58 vdd gnd cell_6t
Xbit_r59_c164 bl_164 br_164 wl_59 vdd gnd cell_6t
Xbit_r60_c164 bl_164 br_164 wl_60 vdd gnd cell_6t
Xbit_r61_c164 bl_164 br_164 wl_61 vdd gnd cell_6t
Xbit_r62_c164 bl_164 br_164 wl_62 vdd gnd cell_6t
Xbit_r63_c164 bl_164 br_164 wl_63 vdd gnd cell_6t
Xbit_r64_c164 bl_164 br_164 wl_64 vdd gnd cell_6t
Xbit_r65_c164 bl_164 br_164 wl_65 vdd gnd cell_6t
Xbit_r66_c164 bl_164 br_164 wl_66 vdd gnd cell_6t
Xbit_r67_c164 bl_164 br_164 wl_67 vdd gnd cell_6t
Xbit_r68_c164 bl_164 br_164 wl_68 vdd gnd cell_6t
Xbit_r69_c164 bl_164 br_164 wl_69 vdd gnd cell_6t
Xbit_r70_c164 bl_164 br_164 wl_70 vdd gnd cell_6t
Xbit_r71_c164 bl_164 br_164 wl_71 vdd gnd cell_6t
Xbit_r72_c164 bl_164 br_164 wl_72 vdd gnd cell_6t
Xbit_r73_c164 bl_164 br_164 wl_73 vdd gnd cell_6t
Xbit_r74_c164 bl_164 br_164 wl_74 vdd gnd cell_6t
Xbit_r75_c164 bl_164 br_164 wl_75 vdd gnd cell_6t
Xbit_r76_c164 bl_164 br_164 wl_76 vdd gnd cell_6t
Xbit_r77_c164 bl_164 br_164 wl_77 vdd gnd cell_6t
Xbit_r78_c164 bl_164 br_164 wl_78 vdd gnd cell_6t
Xbit_r79_c164 bl_164 br_164 wl_79 vdd gnd cell_6t
Xbit_r80_c164 bl_164 br_164 wl_80 vdd gnd cell_6t
Xbit_r81_c164 bl_164 br_164 wl_81 vdd gnd cell_6t
Xbit_r82_c164 bl_164 br_164 wl_82 vdd gnd cell_6t
Xbit_r83_c164 bl_164 br_164 wl_83 vdd gnd cell_6t
Xbit_r84_c164 bl_164 br_164 wl_84 vdd gnd cell_6t
Xbit_r85_c164 bl_164 br_164 wl_85 vdd gnd cell_6t
Xbit_r86_c164 bl_164 br_164 wl_86 vdd gnd cell_6t
Xbit_r87_c164 bl_164 br_164 wl_87 vdd gnd cell_6t
Xbit_r88_c164 bl_164 br_164 wl_88 vdd gnd cell_6t
Xbit_r89_c164 bl_164 br_164 wl_89 vdd gnd cell_6t
Xbit_r90_c164 bl_164 br_164 wl_90 vdd gnd cell_6t
Xbit_r91_c164 bl_164 br_164 wl_91 vdd gnd cell_6t
Xbit_r92_c164 bl_164 br_164 wl_92 vdd gnd cell_6t
Xbit_r93_c164 bl_164 br_164 wl_93 vdd gnd cell_6t
Xbit_r94_c164 bl_164 br_164 wl_94 vdd gnd cell_6t
Xbit_r95_c164 bl_164 br_164 wl_95 vdd gnd cell_6t
Xbit_r96_c164 bl_164 br_164 wl_96 vdd gnd cell_6t
Xbit_r97_c164 bl_164 br_164 wl_97 vdd gnd cell_6t
Xbit_r98_c164 bl_164 br_164 wl_98 vdd gnd cell_6t
Xbit_r99_c164 bl_164 br_164 wl_99 vdd gnd cell_6t
Xbit_r100_c164 bl_164 br_164 wl_100 vdd gnd cell_6t
Xbit_r101_c164 bl_164 br_164 wl_101 vdd gnd cell_6t
Xbit_r102_c164 bl_164 br_164 wl_102 vdd gnd cell_6t
Xbit_r103_c164 bl_164 br_164 wl_103 vdd gnd cell_6t
Xbit_r104_c164 bl_164 br_164 wl_104 vdd gnd cell_6t
Xbit_r105_c164 bl_164 br_164 wl_105 vdd gnd cell_6t
Xbit_r106_c164 bl_164 br_164 wl_106 vdd gnd cell_6t
Xbit_r107_c164 bl_164 br_164 wl_107 vdd gnd cell_6t
Xbit_r108_c164 bl_164 br_164 wl_108 vdd gnd cell_6t
Xbit_r109_c164 bl_164 br_164 wl_109 vdd gnd cell_6t
Xbit_r110_c164 bl_164 br_164 wl_110 vdd gnd cell_6t
Xbit_r111_c164 bl_164 br_164 wl_111 vdd gnd cell_6t
Xbit_r112_c164 bl_164 br_164 wl_112 vdd gnd cell_6t
Xbit_r113_c164 bl_164 br_164 wl_113 vdd gnd cell_6t
Xbit_r114_c164 bl_164 br_164 wl_114 vdd gnd cell_6t
Xbit_r115_c164 bl_164 br_164 wl_115 vdd gnd cell_6t
Xbit_r116_c164 bl_164 br_164 wl_116 vdd gnd cell_6t
Xbit_r117_c164 bl_164 br_164 wl_117 vdd gnd cell_6t
Xbit_r118_c164 bl_164 br_164 wl_118 vdd gnd cell_6t
Xbit_r119_c164 bl_164 br_164 wl_119 vdd gnd cell_6t
Xbit_r120_c164 bl_164 br_164 wl_120 vdd gnd cell_6t
Xbit_r121_c164 bl_164 br_164 wl_121 vdd gnd cell_6t
Xbit_r122_c164 bl_164 br_164 wl_122 vdd gnd cell_6t
Xbit_r123_c164 bl_164 br_164 wl_123 vdd gnd cell_6t
Xbit_r124_c164 bl_164 br_164 wl_124 vdd gnd cell_6t
Xbit_r125_c164 bl_164 br_164 wl_125 vdd gnd cell_6t
Xbit_r126_c164 bl_164 br_164 wl_126 vdd gnd cell_6t
Xbit_r127_c164 bl_164 br_164 wl_127 vdd gnd cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd cell_6t
Xbit_r1_c165 bl_165 br_165 wl_1 vdd gnd cell_6t
Xbit_r2_c165 bl_165 br_165 wl_2 vdd gnd cell_6t
Xbit_r3_c165 bl_165 br_165 wl_3 vdd gnd cell_6t
Xbit_r4_c165 bl_165 br_165 wl_4 vdd gnd cell_6t
Xbit_r5_c165 bl_165 br_165 wl_5 vdd gnd cell_6t
Xbit_r6_c165 bl_165 br_165 wl_6 vdd gnd cell_6t
Xbit_r7_c165 bl_165 br_165 wl_7 vdd gnd cell_6t
Xbit_r8_c165 bl_165 br_165 wl_8 vdd gnd cell_6t
Xbit_r9_c165 bl_165 br_165 wl_9 vdd gnd cell_6t
Xbit_r10_c165 bl_165 br_165 wl_10 vdd gnd cell_6t
Xbit_r11_c165 bl_165 br_165 wl_11 vdd gnd cell_6t
Xbit_r12_c165 bl_165 br_165 wl_12 vdd gnd cell_6t
Xbit_r13_c165 bl_165 br_165 wl_13 vdd gnd cell_6t
Xbit_r14_c165 bl_165 br_165 wl_14 vdd gnd cell_6t
Xbit_r15_c165 bl_165 br_165 wl_15 vdd gnd cell_6t
Xbit_r16_c165 bl_165 br_165 wl_16 vdd gnd cell_6t
Xbit_r17_c165 bl_165 br_165 wl_17 vdd gnd cell_6t
Xbit_r18_c165 bl_165 br_165 wl_18 vdd gnd cell_6t
Xbit_r19_c165 bl_165 br_165 wl_19 vdd gnd cell_6t
Xbit_r20_c165 bl_165 br_165 wl_20 vdd gnd cell_6t
Xbit_r21_c165 bl_165 br_165 wl_21 vdd gnd cell_6t
Xbit_r22_c165 bl_165 br_165 wl_22 vdd gnd cell_6t
Xbit_r23_c165 bl_165 br_165 wl_23 vdd gnd cell_6t
Xbit_r24_c165 bl_165 br_165 wl_24 vdd gnd cell_6t
Xbit_r25_c165 bl_165 br_165 wl_25 vdd gnd cell_6t
Xbit_r26_c165 bl_165 br_165 wl_26 vdd gnd cell_6t
Xbit_r27_c165 bl_165 br_165 wl_27 vdd gnd cell_6t
Xbit_r28_c165 bl_165 br_165 wl_28 vdd gnd cell_6t
Xbit_r29_c165 bl_165 br_165 wl_29 vdd gnd cell_6t
Xbit_r30_c165 bl_165 br_165 wl_30 vdd gnd cell_6t
Xbit_r31_c165 bl_165 br_165 wl_31 vdd gnd cell_6t
Xbit_r32_c165 bl_165 br_165 wl_32 vdd gnd cell_6t
Xbit_r33_c165 bl_165 br_165 wl_33 vdd gnd cell_6t
Xbit_r34_c165 bl_165 br_165 wl_34 vdd gnd cell_6t
Xbit_r35_c165 bl_165 br_165 wl_35 vdd gnd cell_6t
Xbit_r36_c165 bl_165 br_165 wl_36 vdd gnd cell_6t
Xbit_r37_c165 bl_165 br_165 wl_37 vdd gnd cell_6t
Xbit_r38_c165 bl_165 br_165 wl_38 vdd gnd cell_6t
Xbit_r39_c165 bl_165 br_165 wl_39 vdd gnd cell_6t
Xbit_r40_c165 bl_165 br_165 wl_40 vdd gnd cell_6t
Xbit_r41_c165 bl_165 br_165 wl_41 vdd gnd cell_6t
Xbit_r42_c165 bl_165 br_165 wl_42 vdd gnd cell_6t
Xbit_r43_c165 bl_165 br_165 wl_43 vdd gnd cell_6t
Xbit_r44_c165 bl_165 br_165 wl_44 vdd gnd cell_6t
Xbit_r45_c165 bl_165 br_165 wl_45 vdd gnd cell_6t
Xbit_r46_c165 bl_165 br_165 wl_46 vdd gnd cell_6t
Xbit_r47_c165 bl_165 br_165 wl_47 vdd gnd cell_6t
Xbit_r48_c165 bl_165 br_165 wl_48 vdd gnd cell_6t
Xbit_r49_c165 bl_165 br_165 wl_49 vdd gnd cell_6t
Xbit_r50_c165 bl_165 br_165 wl_50 vdd gnd cell_6t
Xbit_r51_c165 bl_165 br_165 wl_51 vdd gnd cell_6t
Xbit_r52_c165 bl_165 br_165 wl_52 vdd gnd cell_6t
Xbit_r53_c165 bl_165 br_165 wl_53 vdd gnd cell_6t
Xbit_r54_c165 bl_165 br_165 wl_54 vdd gnd cell_6t
Xbit_r55_c165 bl_165 br_165 wl_55 vdd gnd cell_6t
Xbit_r56_c165 bl_165 br_165 wl_56 vdd gnd cell_6t
Xbit_r57_c165 bl_165 br_165 wl_57 vdd gnd cell_6t
Xbit_r58_c165 bl_165 br_165 wl_58 vdd gnd cell_6t
Xbit_r59_c165 bl_165 br_165 wl_59 vdd gnd cell_6t
Xbit_r60_c165 bl_165 br_165 wl_60 vdd gnd cell_6t
Xbit_r61_c165 bl_165 br_165 wl_61 vdd gnd cell_6t
Xbit_r62_c165 bl_165 br_165 wl_62 vdd gnd cell_6t
Xbit_r63_c165 bl_165 br_165 wl_63 vdd gnd cell_6t
Xbit_r64_c165 bl_165 br_165 wl_64 vdd gnd cell_6t
Xbit_r65_c165 bl_165 br_165 wl_65 vdd gnd cell_6t
Xbit_r66_c165 bl_165 br_165 wl_66 vdd gnd cell_6t
Xbit_r67_c165 bl_165 br_165 wl_67 vdd gnd cell_6t
Xbit_r68_c165 bl_165 br_165 wl_68 vdd gnd cell_6t
Xbit_r69_c165 bl_165 br_165 wl_69 vdd gnd cell_6t
Xbit_r70_c165 bl_165 br_165 wl_70 vdd gnd cell_6t
Xbit_r71_c165 bl_165 br_165 wl_71 vdd gnd cell_6t
Xbit_r72_c165 bl_165 br_165 wl_72 vdd gnd cell_6t
Xbit_r73_c165 bl_165 br_165 wl_73 vdd gnd cell_6t
Xbit_r74_c165 bl_165 br_165 wl_74 vdd gnd cell_6t
Xbit_r75_c165 bl_165 br_165 wl_75 vdd gnd cell_6t
Xbit_r76_c165 bl_165 br_165 wl_76 vdd gnd cell_6t
Xbit_r77_c165 bl_165 br_165 wl_77 vdd gnd cell_6t
Xbit_r78_c165 bl_165 br_165 wl_78 vdd gnd cell_6t
Xbit_r79_c165 bl_165 br_165 wl_79 vdd gnd cell_6t
Xbit_r80_c165 bl_165 br_165 wl_80 vdd gnd cell_6t
Xbit_r81_c165 bl_165 br_165 wl_81 vdd gnd cell_6t
Xbit_r82_c165 bl_165 br_165 wl_82 vdd gnd cell_6t
Xbit_r83_c165 bl_165 br_165 wl_83 vdd gnd cell_6t
Xbit_r84_c165 bl_165 br_165 wl_84 vdd gnd cell_6t
Xbit_r85_c165 bl_165 br_165 wl_85 vdd gnd cell_6t
Xbit_r86_c165 bl_165 br_165 wl_86 vdd gnd cell_6t
Xbit_r87_c165 bl_165 br_165 wl_87 vdd gnd cell_6t
Xbit_r88_c165 bl_165 br_165 wl_88 vdd gnd cell_6t
Xbit_r89_c165 bl_165 br_165 wl_89 vdd gnd cell_6t
Xbit_r90_c165 bl_165 br_165 wl_90 vdd gnd cell_6t
Xbit_r91_c165 bl_165 br_165 wl_91 vdd gnd cell_6t
Xbit_r92_c165 bl_165 br_165 wl_92 vdd gnd cell_6t
Xbit_r93_c165 bl_165 br_165 wl_93 vdd gnd cell_6t
Xbit_r94_c165 bl_165 br_165 wl_94 vdd gnd cell_6t
Xbit_r95_c165 bl_165 br_165 wl_95 vdd gnd cell_6t
Xbit_r96_c165 bl_165 br_165 wl_96 vdd gnd cell_6t
Xbit_r97_c165 bl_165 br_165 wl_97 vdd gnd cell_6t
Xbit_r98_c165 bl_165 br_165 wl_98 vdd gnd cell_6t
Xbit_r99_c165 bl_165 br_165 wl_99 vdd gnd cell_6t
Xbit_r100_c165 bl_165 br_165 wl_100 vdd gnd cell_6t
Xbit_r101_c165 bl_165 br_165 wl_101 vdd gnd cell_6t
Xbit_r102_c165 bl_165 br_165 wl_102 vdd gnd cell_6t
Xbit_r103_c165 bl_165 br_165 wl_103 vdd gnd cell_6t
Xbit_r104_c165 bl_165 br_165 wl_104 vdd gnd cell_6t
Xbit_r105_c165 bl_165 br_165 wl_105 vdd gnd cell_6t
Xbit_r106_c165 bl_165 br_165 wl_106 vdd gnd cell_6t
Xbit_r107_c165 bl_165 br_165 wl_107 vdd gnd cell_6t
Xbit_r108_c165 bl_165 br_165 wl_108 vdd gnd cell_6t
Xbit_r109_c165 bl_165 br_165 wl_109 vdd gnd cell_6t
Xbit_r110_c165 bl_165 br_165 wl_110 vdd gnd cell_6t
Xbit_r111_c165 bl_165 br_165 wl_111 vdd gnd cell_6t
Xbit_r112_c165 bl_165 br_165 wl_112 vdd gnd cell_6t
Xbit_r113_c165 bl_165 br_165 wl_113 vdd gnd cell_6t
Xbit_r114_c165 bl_165 br_165 wl_114 vdd gnd cell_6t
Xbit_r115_c165 bl_165 br_165 wl_115 vdd gnd cell_6t
Xbit_r116_c165 bl_165 br_165 wl_116 vdd gnd cell_6t
Xbit_r117_c165 bl_165 br_165 wl_117 vdd gnd cell_6t
Xbit_r118_c165 bl_165 br_165 wl_118 vdd gnd cell_6t
Xbit_r119_c165 bl_165 br_165 wl_119 vdd gnd cell_6t
Xbit_r120_c165 bl_165 br_165 wl_120 vdd gnd cell_6t
Xbit_r121_c165 bl_165 br_165 wl_121 vdd gnd cell_6t
Xbit_r122_c165 bl_165 br_165 wl_122 vdd gnd cell_6t
Xbit_r123_c165 bl_165 br_165 wl_123 vdd gnd cell_6t
Xbit_r124_c165 bl_165 br_165 wl_124 vdd gnd cell_6t
Xbit_r125_c165 bl_165 br_165 wl_125 vdd gnd cell_6t
Xbit_r126_c165 bl_165 br_165 wl_126 vdd gnd cell_6t
Xbit_r127_c165 bl_165 br_165 wl_127 vdd gnd cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd cell_6t
Xbit_r1_c166 bl_166 br_166 wl_1 vdd gnd cell_6t
Xbit_r2_c166 bl_166 br_166 wl_2 vdd gnd cell_6t
Xbit_r3_c166 bl_166 br_166 wl_3 vdd gnd cell_6t
Xbit_r4_c166 bl_166 br_166 wl_4 vdd gnd cell_6t
Xbit_r5_c166 bl_166 br_166 wl_5 vdd gnd cell_6t
Xbit_r6_c166 bl_166 br_166 wl_6 vdd gnd cell_6t
Xbit_r7_c166 bl_166 br_166 wl_7 vdd gnd cell_6t
Xbit_r8_c166 bl_166 br_166 wl_8 vdd gnd cell_6t
Xbit_r9_c166 bl_166 br_166 wl_9 vdd gnd cell_6t
Xbit_r10_c166 bl_166 br_166 wl_10 vdd gnd cell_6t
Xbit_r11_c166 bl_166 br_166 wl_11 vdd gnd cell_6t
Xbit_r12_c166 bl_166 br_166 wl_12 vdd gnd cell_6t
Xbit_r13_c166 bl_166 br_166 wl_13 vdd gnd cell_6t
Xbit_r14_c166 bl_166 br_166 wl_14 vdd gnd cell_6t
Xbit_r15_c166 bl_166 br_166 wl_15 vdd gnd cell_6t
Xbit_r16_c166 bl_166 br_166 wl_16 vdd gnd cell_6t
Xbit_r17_c166 bl_166 br_166 wl_17 vdd gnd cell_6t
Xbit_r18_c166 bl_166 br_166 wl_18 vdd gnd cell_6t
Xbit_r19_c166 bl_166 br_166 wl_19 vdd gnd cell_6t
Xbit_r20_c166 bl_166 br_166 wl_20 vdd gnd cell_6t
Xbit_r21_c166 bl_166 br_166 wl_21 vdd gnd cell_6t
Xbit_r22_c166 bl_166 br_166 wl_22 vdd gnd cell_6t
Xbit_r23_c166 bl_166 br_166 wl_23 vdd gnd cell_6t
Xbit_r24_c166 bl_166 br_166 wl_24 vdd gnd cell_6t
Xbit_r25_c166 bl_166 br_166 wl_25 vdd gnd cell_6t
Xbit_r26_c166 bl_166 br_166 wl_26 vdd gnd cell_6t
Xbit_r27_c166 bl_166 br_166 wl_27 vdd gnd cell_6t
Xbit_r28_c166 bl_166 br_166 wl_28 vdd gnd cell_6t
Xbit_r29_c166 bl_166 br_166 wl_29 vdd gnd cell_6t
Xbit_r30_c166 bl_166 br_166 wl_30 vdd gnd cell_6t
Xbit_r31_c166 bl_166 br_166 wl_31 vdd gnd cell_6t
Xbit_r32_c166 bl_166 br_166 wl_32 vdd gnd cell_6t
Xbit_r33_c166 bl_166 br_166 wl_33 vdd gnd cell_6t
Xbit_r34_c166 bl_166 br_166 wl_34 vdd gnd cell_6t
Xbit_r35_c166 bl_166 br_166 wl_35 vdd gnd cell_6t
Xbit_r36_c166 bl_166 br_166 wl_36 vdd gnd cell_6t
Xbit_r37_c166 bl_166 br_166 wl_37 vdd gnd cell_6t
Xbit_r38_c166 bl_166 br_166 wl_38 vdd gnd cell_6t
Xbit_r39_c166 bl_166 br_166 wl_39 vdd gnd cell_6t
Xbit_r40_c166 bl_166 br_166 wl_40 vdd gnd cell_6t
Xbit_r41_c166 bl_166 br_166 wl_41 vdd gnd cell_6t
Xbit_r42_c166 bl_166 br_166 wl_42 vdd gnd cell_6t
Xbit_r43_c166 bl_166 br_166 wl_43 vdd gnd cell_6t
Xbit_r44_c166 bl_166 br_166 wl_44 vdd gnd cell_6t
Xbit_r45_c166 bl_166 br_166 wl_45 vdd gnd cell_6t
Xbit_r46_c166 bl_166 br_166 wl_46 vdd gnd cell_6t
Xbit_r47_c166 bl_166 br_166 wl_47 vdd gnd cell_6t
Xbit_r48_c166 bl_166 br_166 wl_48 vdd gnd cell_6t
Xbit_r49_c166 bl_166 br_166 wl_49 vdd gnd cell_6t
Xbit_r50_c166 bl_166 br_166 wl_50 vdd gnd cell_6t
Xbit_r51_c166 bl_166 br_166 wl_51 vdd gnd cell_6t
Xbit_r52_c166 bl_166 br_166 wl_52 vdd gnd cell_6t
Xbit_r53_c166 bl_166 br_166 wl_53 vdd gnd cell_6t
Xbit_r54_c166 bl_166 br_166 wl_54 vdd gnd cell_6t
Xbit_r55_c166 bl_166 br_166 wl_55 vdd gnd cell_6t
Xbit_r56_c166 bl_166 br_166 wl_56 vdd gnd cell_6t
Xbit_r57_c166 bl_166 br_166 wl_57 vdd gnd cell_6t
Xbit_r58_c166 bl_166 br_166 wl_58 vdd gnd cell_6t
Xbit_r59_c166 bl_166 br_166 wl_59 vdd gnd cell_6t
Xbit_r60_c166 bl_166 br_166 wl_60 vdd gnd cell_6t
Xbit_r61_c166 bl_166 br_166 wl_61 vdd gnd cell_6t
Xbit_r62_c166 bl_166 br_166 wl_62 vdd gnd cell_6t
Xbit_r63_c166 bl_166 br_166 wl_63 vdd gnd cell_6t
Xbit_r64_c166 bl_166 br_166 wl_64 vdd gnd cell_6t
Xbit_r65_c166 bl_166 br_166 wl_65 vdd gnd cell_6t
Xbit_r66_c166 bl_166 br_166 wl_66 vdd gnd cell_6t
Xbit_r67_c166 bl_166 br_166 wl_67 vdd gnd cell_6t
Xbit_r68_c166 bl_166 br_166 wl_68 vdd gnd cell_6t
Xbit_r69_c166 bl_166 br_166 wl_69 vdd gnd cell_6t
Xbit_r70_c166 bl_166 br_166 wl_70 vdd gnd cell_6t
Xbit_r71_c166 bl_166 br_166 wl_71 vdd gnd cell_6t
Xbit_r72_c166 bl_166 br_166 wl_72 vdd gnd cell_6t
Xbit_r73_c166 bl_166 br_166 wl_73 vdd gnd cell_6t
Xbit_r74_c166 bl_166 br_166 wl_74 vdd gnd cell_6t
Xbit_r75_c166 bl_166 br_166 wl_75 vdd gnd cell_6t
Xbit_r76_c166 bl_166 br_166 wl_76 vdd gnd cell_6t
Xbit_r77_c166 bl_166 br_166 wl_77 vdd gnd cell_6t
Xbit_r78_c166 bl_166 br_166 wl_78 vdd gnd cell_6t
Xbit_r79_c166 bl_166 br_166 wl_79 vdd gnd cell_6t
Xbit_r80_c166 bl_166 br_166 wl_80 vdd gnd cell_6t
Xbit_r81_c166 bl_166 br_166 wl_81 vdd gnd cell_6t
Xbit_r82_c166 bl_166 br_166 wl_82 vdd gnd cell_6t
Xbit_r83_c166 bl_166 br_166 wl_83 vdd gnd cell_6t
Xbit_r84_c166 bl_166 br_166 wl_84 vdd gnd cell_6t
Xbit_r85_c166 bl_166 br_166 wl_85 vdd gnd cell_6t
Xbit_r86_c166 bl_166 br_166 wl_86 vdd gnd cell_6t
Xbit_r87_c166 bl_166 br_166 wl_87 vdd gnd cell_6t
Xbit_r88_c166 bl_166 br_166 wl_88 vdd gnd cell_6t
Xbit_r89_c166 bl_166 br_166 wl_89 vdd gnd cell_6t
Xbit_r90_c166 bl_166 br_166 wl_90 vdd gnd cell_6t
Xbit_r91_c166 bl_166 br_166 wl_91 vdd gnd cell_6t
Xbit_r92_c166 bl_166 br_166 wl_92 vdd gnd cell_6t
Xbit_r93_c166 bl_166 br_166 wl_93 vdd gnd cell_6t
Xbit_r94_c166 bl_166 br_166 wl_94 vdd gnd cell_6t
Xbit_r95_c166 bl_166 br_166 wl_95 vdd gnd cell_6t
Xbit_r96_c166 bl_166 br_166 wl_96 vdd gnd cell_6t
Xbit_r97_c166 bl_166 br_166 wl_97 vdd gnd cell_6t
Xbit_r98_c166 bl_166 br_166 wl_98 vdd gnd cell_6t
Xbit_r99_c166 bl_166 br_166 wl_99 vdd gnd cell_6t
Xbit_r100_c166 bl_166 br_166 wl_100 vdd gnd cell_6t
Xbit_r101_c166 bl_166 br_166 wl_101 vdd gnd cell_6t
Xbit_r102_c166 bl_166 br_166 wl_102 vdd gnd cell_6t
Xbit_r103_c166 bl_166 br_166 wl_103 vdd gnd cell_6t
Xbit_r104_c166 bl_166 br_166 wl_104 vdd gnd cell_6t
Xbit_r105_c166 bl_166 br_166 wl_105 vdd gnd cell_6t
Xbit_r106_c166 bl_166 br_166 wl_106 vdd gnd cell_6t
Xbit_r107_c166 bl_166 br_166 wl_107 vdd gnd cell_6t
Xbit_r108_c166 bl_166 br_166 wl_108 vdd gnd cell_6t
Xbit_r109_c166 bl_166 br_166 wl_109 vdd gnd cell_6t
Xbit_r110_c166 bl_166 br_166 wl_110 vdd gnd cell_6t
Xbit_r111_c166 bl_166 br_166 wl_111 vdd gnd cell_6t
Xbit_r112_c166 bl_166 br_166 wl_112 vdd gnd cell_6t
Xbit_r113_c166 bl_166 br_166 wl_113 vdd gnd cell_6t
Xbit_r114_c166 bl_166 br_166 wl_114 vdd gnd cell_6t
Xbit_r115_c166 bl_166 br_166 wl_115 vdd gnd cell_6t
Xbit_r116_c166 bl_166 br_166 wl_116 vdd gnd cell_6t
Xbit_r117_c166 bl_166 br_166 wl_117 vdd gnd cell_6t
Xbit_r118_c166 bl_166 br_166 wl_118 vdd gnd cell_6t
Xbit_r119_c166 bl_166 br_166 wl_119 vdd gnd cell_6t
Xbit_r120_c166 bl_166 br_166 wl_120 vdd gnd cell_6t
Xbit_r121_c166 bl_166 br_166 wl_121 vdd gnd cell_6t
Xbit_r122_c166 bl_166 br_166 wl_122 vdd gnd cell_6t
Xbit_r123_c166 bl_166 br_166 wl_123 vdd gnd cell_6t
Xbit_r124_c166 bl_166 br_166 wl_124 vdd gnd cell_6t
Xbit_r125_c166 bl_166 br_166 wl_125 vdd gnd cell_6t
Xbit_r126_c166 bl_166 br_166 wl_126 vdd gnd cell_6t
Xbit_r127_c166 bl_166 br_166 wl_127 vdd gnd cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd cell_6t
Xbit_r1_c167 bl_167 br_167 wl_1 vdd gnd cell_6t
Xbit_r2_c167 bl_167 br_167 wl_2 vdd gnd cell_6t
Xbit_r3_c167 bl_167 br_167 wl_3 vdd gnd cell_6t
Xbit_r4_c167 bl_167 br_167 wl_4 vdd gnd cell_6t
Xbit_r5_c167 bl_167 br_167 wl_5 vdd gnd cell_6t
Xbit_r6_c167 bl_167 br_167 wl_6 vdd gnd cell_6t
Xbit_r7_c167 bl_167 br_167 wl_7 vdd gnd cell_6t
Xbit_r8_c167 bl_167 br_167 wl_8 vdd gnd cell_6t
Xbit_r9_c167 bl_167 br_167 wl_9 vdd gnd cell_6t
Xbit_r10_c167 bl_167 br_167 wl_10 vdd gnd cell_6t
Xbit_r11_c167 bl_167 br_167 wl_11 vdd gnd cell_6t
Xbit_r12_c167 bl_167 br_167 wl_12 vdd gnd cell_6t
Xbit_r13_c167 bl_167 br_167 wl_13 vdd gnd cell_6t
Xbit_r14_c167 bl_167 br_167 wl_14 vdd gnd cell_6t
Xbit_r15_c167 bl_167 br_167 wl_15 vdd gnd cell_6t
Xbit_r16_c167 bl_167 br_167 wl_16 vdd gnd cell_6t
Xbit_r17_c167 bl_167 br_167 wl_17 vdd gnd cell_6t
Xbit_r18_c167 bl_167 br_167 wl_18 vdd gnd cell_6t
Xbit_r19_c167 bl_167 br_167 wl_19 vdd gnd cell_6t
Xbit_r20_c167 bl_167 br_167 wl_20 vdd gnd cell_6t
Xbit_r21_c167 bl_167 br_167 wl_21 vdd gnd cell_6t
Xbit_r22_c167 bl_167 br_167 wl_22 vdd gnd cell_6t
Xbit_r23_c167 bl_167 br_167 wl_23 vdd gnd cell_6t
Xbit_r24_c167 bl_167 br_167 wl_24 vdd gnd cell_6t
Xbit_r25_c167 bl_167 br_167 wl_25 vdd gnd cell_6t
Xbit_r26_c167 bl_167 br_167 wl_26 vdd gnd cell_6t
Xbit_r27_c167 bl_167 br_167 wl_27 vdd gnd cell_6t
Xbit_r28_c167 bl_167 br_167 wl_28 vdd gnd cell_6t
Xbit_r29_c167 bl_167 br_167 wl_29 vdd gnd cell_6t
Xbit_r30_c167 bl_167 br_167 wl_30 vdd gnd cell_6t
Xbit_r31_c167 bl_167 br_167 wl_31 vdd gnd cell_6t
Xbit_r32_c167 bl_167 br_167 wl_32 vdd gnd cell_6t
Xbit_r33_c167 bl_167 br_167 wl_33 vdd gnd cell_6t
Xbit_r34_c167 bl_167 br_167 wl_34 vdd gnd cell_6t
Xbit_r35_c167 bl_167 br_167 wl_35 vdd gnd cell_6t
Xbit_r36_c167 bl_167 br_167 wl_36 vdd gnd cell_6t
Xbit_r37_c167 bl_167 br_167 wl_37 vdd gnd cell_6t
Xbit_r38_c167 bl_167 br_167 wl_38 vdd gnd cell_6t
Xbit_r39_c167 bl_167 br_167 wl_39 vdd gnd cell_6t
Xbit_r40_c167 bl_167 br_167 wl_40 vdd gnd cell_6t
Xbit_r41_c167 bl_167 br_167 wl_41 vdd gnd cell_6t
Xbit_r42_c167 bl_167 br_167 wl_42 vdd gnd cell_6t
Xbit_r43_c167 bl_167 br_167 wl_43 vdd gnd cell_6t
Xbit_r44_c167 bl_167 br_167 wl_44 vdd gnd cell_6t
Xbit_r45_c167 bl_167 br_167 wl_45 vdd gnd cell_6t
Xbit_r46_c167 bl_167 br_167 wl_46 vdd gnd cell_6t
Xbit_r47_c167 bl_167 br_167 wl_47 vdd gnd cell_6t
Xbit_r48_c167 bl_167 br_167 wl_48 vdd gnd cell_6t
Xbit_r49_c167 bl_167 br_167 wl_49 vdd gnd cell_6t
Xbit_r50_c167 bl_167 br_167 wl_50 vdd gnd cell_6t
Xbit_r51_c167 bl_167 br_167 wl_51 vdd gnd cell_6t
Xbit_r52_c167 bl_167 br_167 wl_52 vdd gnd cell_6t
Xbit_r53_c167 bl_167 br_167 wl_53 vdd gnd cell_6t
Xbit_r54_c167 bl_167 br_167 wl_54 vdd gnd cell_6t
Xbit_r55_c167 bl_167 br_167 wl_55 vdd gnd cell_6t
Xbit_r56_c167 bl_167 br_167 wl_56 vdd gnd cell_6t
Xbit_r57_c167 bl_167 br_167 wl_57 vdd gnd cell_6t
Xbit_r58_c167 bl_167 br_167 wl_58 vdd gnd cell_6t
Xbit_r59_c167 bl_167 br_167 wl_59 vdd gnd cell_6t
Xbit_r60_c167 bl_167 br_167 wl_60 vdd gnd cell_6t
Xbit_r61_c167 bl_167 br_167 wl_61 vdd gnd cell_6t
Xbit_r62_c167 bl_167 br_167 wl_62 vdd gnd cell_6t
Xbit_r63_c167 bl_167 br_167 wl_63 vdd gnd cell_6t
Xbit_r64_c167 bl_167 br_167 wl_64 vdd gnd cell_6t
Xbit_r65_c167 bl_167 br_167 wl_65 vdd gnd cell_6t
Xbit_r66_c167 bl_167 br_167 wl_66 vdd gnd cell_6t
Xbit_r67_c167 bl_167 br_167 wl_67 vdd gnd cell_6t
Xbit_r68_c167 bl_167 br_167 wl_68 vdd gnd cell_6t
Xbit_r69_c167 bl_167 br_167 wl_69 vdd gnd cell_6t
Xbit_r70_c167 bl_167 br_167 wl_70 vdd gnd cell_6t
Xbit_r71_c167 bl_167 br_167 wl_71 vdd gnd cell_6t
Xbit_r72_c167 bl_167 br_167 wl_72 vdd gnd cell_6t
Xbit_r73_c167 bl_167 br_167 wl_73 vdd gnd cell_6t
Xbit_r74_c167 bl_167 br_167 wl_74 vdd gnd cell_6t
Xbit_r75_c167 bl_167 br_167 wl_75 vdd gnd cell_6t
Xbit_r76_c167 bl_167 br_167 wl_76 vdd gnd cell_6t
Xbit_r77_c167 bl_167 br_167 wl_77 vdd gnd cell_6t
Xbit_r78_c167 bl_167 br_167 wl_78 vdd gnd cell_6t
Xbit_r79_c167 bl_167 br_167 wl_79 vdd gnd cell_6t
Xbit_r80_c167 bl_167 br_167 wl_80 vdd gnd cell_6t
Xbit_r81_c167 bl_167 br_167 wl_81 vdd gnd cell_6t
Xbit_r82_c167 bl_167 br_167 wl_82 vdd gnd cell_6t
Xbit_r83_c167 bl_167 br_167 wl_83 vdd gnd cell_6t
Xbit_r84_c167 bl_167 br_167 wl_84 vdd gnd cell_6t
Xbit_r85_c167 bl_167 br_167 wl_85 vdd gnd cell_6t
Xbit_r86_c167 bl_167 br_167 wl_86 vdd gnd cell_6t
Xbit_r87_c167 bl_167 br_167 wl_87 vdd gnd cell_6t
Xbit_r88_c167 bl_167 br_167 wl_88 vdd gnd cell_6t
Xbit_r89_c167 bl_167 br_167 wl_89 vdd gnd cell_6t
Xbit_r90_c167 bl_167 br_167 wl_90 vdd gnd cell_6t
Xbit_r91_c167 bl_167 br_167 wl_91 vdd gnd cell_6t
Xbit_r92_c167 bl_167 br_167 wl_92 vdd gnd cell_6t
Xbit_r93_c167 bl_167 br_167 wl_93 vdd gnd cell_6t
Xbit_r94_c167 bl_167 br_167 wl_94 vdd gnd cell_6t
Xbit_r95_c167 bl_167 br_167 wl_95 vdd gnd cell_6t
Xbit_r96_c167 bl_167 br_167 wl_96 vdd gnd cell_6t
Xbit_r97_c167 bl_167 br_167 wl_97 vdd gnd cell_6t
Xbit_r98_c167 bl_167 br_167 wl_98 vdd gnd cell_6t
Xbit_r99_c167 bl_167 br_167 wl_99 vdd gnd cell_6t
Xbit_r100_c167 bl_167 br_167 wl_100 vdd gnd cell_6t
Xbit_r101_c167 bl_167 br_167 wl_101 vdd gnd cell_6t
Xbit_r102_c167 bl_167 br_167 wl_102 vdd gnd cell_6t
Xbit_r103_c167 bl_167 br_167 wl_103 vdd gnd cell_6t
Xbit_r104_c167 bl_167 br_167 wl_104 vdd gnd cell_6t
Xbit_r105_c167 bl_167 br_167 wl_105 vdd gnd cell_6t
Xbit_r106_c167 bl_167 br_167 wl_106 vdd gnd cell_6t
Xbit_r107_c167 bl_167 br_167 wl_107 vdd gnd cell_6t
Xbit_r108_c167 bl_167 br_167 wl_108 vdd gnd cell_6t
Xbit_r109_c167 bl_167 br_167 wl_109 vdd gnd cell_6t
Xbit_r110_c167 bl_167 br_167 wl_110 vdd gnd cell_6t
Xbit_r111_c167 bl_167 br_167 wl_111 vdd gnd cell_6t
Xbit_r112_c167 bl_167 br_167 wl_112 vdd gnd cell_6t
Xbit_r113_c167 bl_167 br_167 wl_113 vdd gnd cell_6t
Xbit_r114_c167 bl_167 br_167 wl_114 vdd gnd cell_6t
Xbit_r115_c167 bl_167 br_167 wl_115 vdd gnd cell_6t
Xbit_r116_c167 bl_167 br_167 wl_116 vdd gnd cell_6t
Xbit_r117_c167 bl_167 br_167 wl_117 vdd gnd cell_6t
Xbit_r118_c167 bl_167 br_167 wl_118 vdd gnd cell_6t
Xbit_r119_c167 bl_167 br_167 wl_119 vdd gnd cell_6t
Xbit_r120_c167 bl_167 br_167 wl_120 vdd gnd cell_6t
Xbit_r121_c167 bl_167 br_167 wl_121 vdd gnd cell_6t
Xbit_r122_c167 bl_167 br_167 wl_122 vdd gnd cell_6t
Xbit_r123_c167 bl_167 br_167 wl_123 vdd gnd cell_6t
Xbit_r124_c167 bl_167 br_167 wl_124 vdd gnd cell_6t
Xbit_r125_c167 bl_167 br_167 wl_125 vdd gnd cell_6t
Xbit_r126_c167 bl_167 br_167 wl_126 vdd gnd cell_6t
Xbit_r127_c167 bl_167 br_167 wl_127 vdd gnd cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd cell_6t
Xbit_r1_c168 bl_168 br_168 wl_1 vdd gnd cell_6t
Xbit_r2_c168 bl_168 br_168 wl_2 vdd gnd cell_6t
Xbit_r3_c168 bl_168 br_168 wl_3 vdd gnd cell_6t
Xbit_r4_c168 bl_168 br_168 wl_4 vdd gnd cell_6t
Xbit_r5_c168 bl_168 br_168 wl_5 vdd gnd cell_6t
Xbit_r6_c168 bl_168 br_168 wl_6 vdd gnd cell_6t
Xbit_r7_c168 bl_168 br_168 wl_7 vdd gnd cell_6t
Xbit_r8_c168 bl_168 br_168 wl_8 vdd gnd cell_6t
Xbit_r9_c168 bl_168 br_168 wl_9 vdd gnd cell_6t
Xbit_r10_c168 bl_168 br_168 wl_10 vdd gnd cell_6t
Xbit_r11_c168 bl_168 br_168 wl_11 vdd gnd cell_6t
Xbit_r12_c168 bl_168 br_168 wl_12 vdd gnd cell_6t
Xbit_r13_c168 bl_168 br_168 wl_13 vdd gnd cell_6t
Xbit_r14_c168 bl_168 br_168 wl_14 vdd gnd cell_6t
Xbit_r15_c168 bl_168 br_168 wl_15 vdd gnd cell_6t
Xbit_r16_c168 bl_168 br_168 wl_16 vdd gnd cell_6t
Xbit_r17_c168 bl_168 br_168 wl_17 vdd gnd cell_6t
Xbit_r18_c168 bl_168 br_168 wl_18 vdd gnd cell_6t
Xbit_r19_c168 bl_168 br_168 wl_19 vdd gnd cell_6t
Xbit_r20_c168 bl_168 br_168 wl_20 vdd gnd cell_6t
Xbit_r21_c168 bl_168 br_168 wl_21 vdd gnd cell_6t
Xbit_r22_c168 bl_168 br_168 wl_22 vdd gnd cell_6t
Xbit_r23_c168 bl_168 br_168 wl_23 vdd gnd cell_6t
Xbit_r24_c168 bl_168 br_168 wl_24 vdd gnd cell_6t
Xbit_r25_c168 bl_168 br_168 wl_25 vdd gnd cell_6t
Xbit_r26_c168 bl_168 br_168 wl_26 vdd gnd cell_6t
Xbit_r27_c168 bl_168 br_168 wl_27 vdd gnd cell_6t
Xbit_r28_c168 bl_168 br_168 wl_28 vdd gnd cell_6t
Xbit_r29_c168 bl_168 br_168 wl_29 vdd gnd cell_6t
Xbit_r30_c168 bl_168 br_168 wl_30 vdd gnd cell_6t
Xbit_r31_c168 bl_168 br_168 wl_31 vdd gnd cell_6t
Xbit_r32_c168 bl_168 br_168 wl_32 vdd gnd cell_6t
Xbit_r33_c168 bl_168 br_168 wl_33 vdd gnd cell_6t
Xbit_r34_c168 bl_168 br_168 wl_34 vdd gnd cell_6t
Xbit_r35_c168 bl_168 br_168 wl_35 vdd gnd cell_6t
Xbit_r36_c168 bl_168 br_168 wl_36 vdd gnd cell_6t
Xbit_r37_c168 bl_168 br_168 wl_37 vdd gnd cell_6t
Xbit_r38_c168 bl_168 br_168 wl_38 vdd gnd cell_6t
Xbit_r39_c168 bl_168 br_168 wl_39 vdd gnd cell_6t
Xbit_r40_c168 bl_168 br_168 wl_40 vdd gnd cell_6t
Xbit_r41_c168 bl_168 br_168 wl_41 vdd gnd cell_6t
Xbit_r42_c168 bl_168 br_168 wl_42 vdd gnd cell_6t
Xbit_r43_c168 bl_168 br_168 wl_43 vdd gnd cell_6t
Xbit_r44_c168 bl_168 br_168 wl_44 vdd gnd cell_6t
Xbit_r45_c168 bl_168 br_168 wl_45 vdd gnd cell_6t
Xbit_r46_c168 bl_168 br_168 wl_46 vdd gnd cell_6t
Xbit_r47_c168 bl_168 br_168 wl_47 vdd gnd cell_6t
Xbit_r48_c168 bl_168 br_168 wl_48 vdd gnd cell_6t
Xbit_r49_c168 bl_168 br_168 wl_49 vdd gnd cell_6t
Xbit_r50_c168 bl_168 br_168 wl_50 vdd gnd cell_6t
Xbit_r51_c168 bl_168 br_168 wl_51 vdd gnd cell_6t
Xbit_r52_c168 bl_168 br_168 wl_52 vdd gnd cell_6t
Xbit_r53_c168 bl_168 br_168 wl_53 vdd gnd cell_6t
Xbit_r54_c168 bl_168 br_168 wl_54 vdd gnd cell_6t
Xbit_r55_c168 bl_168 br_168 wl_55 vdd gnd cell_6t
Xbit_r56_c168 bl_168 br_168 wl_56 vdd gnd cell_6t
Xbit_r57_c168 bl_168 br_168 wl_57 vdd gnd cell_6t
Xbit_r58_c168 bl_168 br_168 wl_58 vdd gnd cell_6t
Xbit_r59_c168 bl_168 br_168 wl_59 vdd gnd cell_6t
Xbit_r60_c168 bl_168 br_168 wl_60 vdd gnd cell_6t
Xbit_r61_c168 bl_168 br_168 wl_61 vdd gnd cell_6t
Xbit_r62_c168 bl_168 br_168 wl_62 vdd gnd cell_6t
Xbit_r63_c168 bl_168 br_168 wl_63 vdd gnd cell_6t
Xbit_r64_c168 bl_168 br_168 wl_64 vdd gnd cell_6t
Xbit_r65_c168 bl_168 br_168 wl_65 vdd gnd cell_6t
Xbit_r66_c168 bl_168 br_168 wl_66 vdd gnd cell_6t
Xbit_r67_c168 bl_168 br_168 wl_67 vdd gnd cell_6t
Xbit_r68_c168 bl_168 br_168 wl_68 vdd gnd cell_6t
Xbit_r69_c168 bl_168 br_168 wl_69 vdd gnd cell_6t
Xbit_r70_c168 bl_168 br_168 wl_70 vdd gnd cell_6t
Xbit_r71_c168 bl_168 br_168 wl_71 vdd gnd cell_6t
Xbit_r72_c168 bl_168 br_168 wl_72 vdd gnd cell_6t
Xbit_r73_c168 bl_168 br_168 wl_73 vdd gnd cell_6t
Xbit_r74_c168 bl_168 br_168 wl_74 vdd gnd cell_6t
Xbit_r75_c168 bl_168 br_168 wl_75 vdd gnd cell_6t
Xbit_r76_c168 bl_168 br_168 wl_76 vdd gnd cell_6t
Xbit_r77_c168 bl_168 br_168 wl_77 vdd gnd cell_6t
Xbit_r78_c168 bl_168 br_168 wl_78 vdd gnd cell_6t
Xbit_r79_c168 bl_168 br_168 wl_79 vdd gnd cell_6t
Xbit_r80_c168 bl_168 br_168 wl_80 vdd gnd cell_6t
Xbit_r81_c168 bl_168 br_168 wl_81 vdd gnd cell_6t
Xbit_r82_c168 bl_168 br_168 wl_82 vdd gnd cell_6t
Xbit_r83_c168 bl_168 br_168 wl_83 vdd gnd cell_6t
Xbit_r84_c168 bl_168 br_168 wl_84 vdd gnd cell_6t
Xbit_r85_c168 bl_168 br_168 wl_85 vdd gnd cell_6t
Xbit_r86_c168 bl_168 br_168 wl_86 vdd gnd cell_6t
Xbit_r87_c168 bl_168 br_168 wl_87 vdd gnd cell_6t
Xbit_r88_c168 bl_168 br_168 wl_88 vdd gnd cell_6t
Xbit_r89_c168 bl_168 br_168 wl_89 vdd gnd cell_6t
Xbit_r90_c168 bl_168 br_168 wl_90 vdd gnd cell_6t
Xbit_r91_c168 bl_168 br_168 wl_91 vdd gnd cell_6t
Xbit_r92_c168 bl_168 br_168 wl_92 vdd gnd cell_6t
Xbit_r93_c168 bl_168 br_168 wl_93 vdd gnd cell_6t
Xbit_r94_c168 bl_168 br_168 wl_94 vdd gnd cell_6t
Xbit_r95_c168 bl_168 br_168 wl_95 vdd gnd cell_6t
Xbit_r96_c168 bl_168 br_168 wl_96 vdd gnd cell_6t
Xbit_r97_c168 bl_168 br_168 wl_97 vdd gnd cell_6t
Xbit_r98_c168 bl_168 br_168 wl_98 vdd gnd cell_6t
Xbit_r99_c168 bl_168 br_168 wl_99 vdd gnd cell_6t
Xbit_r100_c168 bl_168 br_168 wl_100 vdd gnd cell_6t
Xbit_r101_c168 bl_168 br_168 wl_101 vdd gnd cell_6t
Xbit_r102_c168 bl_168 br_168 wl_102 vdd gnd cell_6t
Xbit_r103_c168 bl_168 br_168 wl_103 vdd gnd cell_6t
Xbit_r104_c168 bl_168 br_168 wl_104 vdd gnd cell_6t
Xbit_r105_c168 bl_168 br_168 wl_105 vdd gnd cell_6t
Xbit_r106_c168 bl_168 br_168 wl_106 vdd gnd cell_6t
Xbit_r107_c168 bl_168 br_168 wl_107 vdd gnd cell_6t
Xbit_r108_c168 bl_168 br_168 wl_108 vdd gnd cell_6t
Xbit_r109_c168 bl_168 br_168 wl_109 vdd gnd cell_6t
Xbit_r110_c168 bl_168 br_168 wl_110 vdd gnd cell_6t
Xbit_r111_c168 bl_168 br_168 wl_111 vdd gnd cell_6t
Xbit_r112_c168 bl_168 br_168 wl_112 vdd gnd cell_6t
Xbit_r113_c168 bl_168 br_168 wl_113 vdd gnd cell_6t
Xbit_r114_c168 bl_168 br_168 wl_114 vdd gnd cell_6t
Xbit_r115_c168 bl_168 br_168 wl_115 vdd gnd cell_6t
Xbit_r116_c168 bl_168 br_168 wl_116 vdd gnd cell_6t
Xbit_r117_c168 bl_168 br_168 wl_117 vdd gnd cell_6t
Xbit_r118_c168 bl_168 br_168 wl_118 vdd gnd cell_6t
Xbit_r119_c168 bl_168 br_168 wl_119 vdd gnd cell_6t
Xbit_r120_c168 bl_168 br_168 wl_120 vdd gnd cell_6t
Xbit_r121_c168 bl_168 br_168 wl_121 vdd gnd cell_6t
Xbit_r122_c168 bl_168 br_168 wl_122 vdd gnd cell_6t
Xbit_r123_c168 bl_168 br_168 wl_123 vdd gnd cell_6t
Xbit_r124_c168 bl_168 br_168 wl_124 vdd gnd cell_6t
Xbit_r125_c168 bl_168 br_168 wl_125 vdd gnd cell_6t
Xbit_r126_c168 bl_168 br_168 wl_126 vdd gnd cell_6t
Xbit_r127_c168 bl_168 br_168 wl_127 vdd gnd cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd cell_6t
Xbit_r1_c169 bl_169 br_169 wl_1 vdd gnd cell_6t
Xbit_r2_c169 bl_169 br_169 wl_2 vdd gnd cell_6t
Xbit_r3_c169 bl_169 br_169 wl_3 vdd gnd cell_6t
Xbit_r4_c169 bl_169 br_169 wl_4 vdd gnd cell_6t
Xbit_r5_c169 bl_169 br_169 wl_5 vdd gnd cell_6t
Xbit_r6_c169 bl_169 br_169 wl_6 vdd gnd cell_6t
Xbit_r7_c169 bl_169 br_169 wl_7 vdd gnd cell_6t
Xbit_r8_c169 bl_169 br_169 wl_8 vdd gnd cell_6t
Xbit_r9_c169 bl_169 br_169 wl_9 vdd gnd cell_6t
Xbit_r10_c169 bl_169 br_169 wl_10 vdd gnd cell_6t
Xbit_r11_c169 bl_169 br_169 wl_11 vdd gnd cell_6t
Xbit_r12_c169 bl_169 br_169 wl_12 vdd gnd cell_6t
Xbit_r13_c169 bl_169 br_169 wl_13 vdd gnd cell_6t
Xbit_r14_c169 bl_169 br_169 wl_14 vdd gnd cell_6t
Xbit_r15_c169 bl_169 br_169 wl_15 vdd gnd cell_6t
Xbit_r16_c169 bl_169 br_169 wl_16 vdd gnd cell_6t
Xbit_r17_c169 bl_169 br_169 wl_17 vdd gnd cell_6t
Xbit_r18_c169 bl_169 br_169 wl_18 vdd gnd cell_6t
Xbit_r19_c169 bl_169 br_169 wl_19 vdd gnd cell_6t
Xbit_r20_c169 bl_169 br_169 wl_20 vdd gnd cell_6t
Xbit_r21_c169 bl_169 br_169 wl_21 vdd gnd cell_6t
Xbit_r22_c169 bl_169 br_169 wl_22 vdd gnd cell_6t
Xbit_r23_c169 bl_169 br_169 wl_23 vdd gnd cell_6t
Xbit_r24_c169 bl_169 br_169 wl_24 vdd gnd cell_6t
Xbit_r25_c169 bl_169 br_169 wl_25 vdd gnd cell_6t
Xbit_r26_c169 bl_169 br_169 wl_26 vdd gnd cell_6t
Xbit_r27_c169 bl_169 br_169 wl_27 vdd gnd cell_6t
Xbit_r28_c169 bl_169 br_169 wl_28 vdd gnd cell_6t
Xbit_r29_c169 bl_169 br_169 wl_29 vdd gnd cell_6t
Xbit_r30_c169 bl_169 br_169 wl_30 vdd gnd cell_6t
Xbit_r31_c169 bl_169 br_169 wl_31 vdd gnd cell_6t
Xbit_r32_c169 bl_169 br_169 wl_32 vdd gnd cell_6t
Xbit_r33_c169 bl_169 br_169 wl_33 vdd gnd cell_6t
Xbit_r34_c169 bl_169 br_169 wl_34 vdd gnd cell_6t
Xbit_r35_c169 bl_169 br_169 wl_35 vdd gnd cell_6t
Xbit_r36_c169 bl_169 br_169 wl_36 vdd gnd cell_6t
Xbit_r37_c169 bl_169 br_169 wl_37 vdd gnd cell_6t
Xbit_r38_c169 bl_169 br_169 wl_38 vdd gnd cell_6t
Xbit_r39_c169 bl_169 br_169 wl_39 vdd gnd cell_6t
Xbit_r40_c169 bl_169 br_169 wl_40 vdd gnd cell_6t
Xbit_r41_c169 bl_169 br_169 wl_41 vdd gnd cell_6t
Xbit_r42_c169 bl_169 br_169 wl_42 vdd gnd cell_6t
Xbit_r43_c169 bl_169 br_169 wl_43 vdd gnd cell_6t
Xbit_r44_c169 bl_169 br_169 wl_44 vdd gnd cell_6t
Xbit_r45_c169 bl_169 br_169 wl_45 vdd gnd cell_6t
Xbit_r46_c169 bl_169 br_169 wl_46 vdd gnd cell_6t
Xbit_r47_c169 bl_169 br_169 wl_47 vdd gnd cell_6t
Xbit_r48_c169 bl_169 br_169 wl_48 vdd gnd cell_6t
Xbit_r49_c169 bl_169 br_169 wl_49 vdd gnd cell_6t
Xbit_r50_c169 bl_169 br_169 wl_50 vdd gnd cell_6t
Xbit_r51_c169 bl_169 br_169 wl_51 vdd gnd cell_6t
Xbit_r52_c169 bl_169 br_169 wl_52 vdd gnd cell_6t
Xbit_r53_c169 bl_169 br_169 wl_53 vdd gnd cell_6t
Xbit_r54_c169 bl_169 br_169 wl_54 vdd gnd cell_6t
Xbit_r55_c169 bl_169 br_169 wl_55 vdd gnd cell_6t
Xbit_r56_c169 bl_169 br_169 wl_56 vdd gnd cell_6t
Xbit_r57_c169 bl_169 br_169 wl_57 vdd gnd cell_6t
Xbit_r58_c169 bl_169 br_169 wl_58 vdd gnd cell_6t
Xbit_r59_c169 bl_169 br_169 wl_59 vdd gnd cell_6t
Xbit_r60_c169 bl_169 br_169 wl_60 vdd gnd cell_6t
Xbit_r61_c169 bl_169 br_169 wl_61 vdd gnd cell_6t
Xbit_r62_c169 bl_169 br_169 wl_62 vdd gnd cell_6t
Xbit_r63_c169 bl_169 br_169 wl_63 vdd gnd cell_6t
Xbit_r64_c169 bl_169 br_169 wl_64 vdd gnd cell_6t
Xbit_r65_c169 bl_169 br_169 wl_65 vdd gnd cell_6t
Xbit_r66_c169 bl_169 br_169 wl_66 vdd gnd cell_6t
Xbit_r67_c169 bl_169 br_169 wl_67 vdd gnd cell_6t
Xbit_r68_c169 bl_169 br_169 wl_68 vdd gnd cell_6t
Xbit_r69_c169 bl_169 br_169 wl_69 vdd gnd cell_6t
Xbit_r70_c169 bl_169 br_169 wl_70 vdd gnd cell_6t
Xbit_r71_c169 bl_169 br_169 wl_71 vdd gnd cell_6t
Xbit_r72_c169 bl_169 br_169 wl_72 vdd gnd cell_6t
Xbit_r73_c169 bl_169 br_169 wl_73 vdd gnd cell_6t
Xbit_r74_c169 bl_169 br_169 wl_74 vdd gnd cell_6t
Xbit_r75_c169 bl_169 br_169 wl_75 vdd gnd cell_6t
Xbit_r76_c169 bl_169 br_169 wl_76 vdd gnd cell_6t
Xbit_r77_c169 bl_169 br_169 wl_77 vdd gnd cell_6t
Xbit_r78_c169 bl_169 br_169 wl_78 vdd gnd cell_6t
Xbit_r79_c169 bl_169 br_169 wl_79 vdd gnd cell_6t
Xbit_r80_c169 bl_169 br_169 wl_80 vdd gnd cell_6t
Xbit_r81_c169 bl_169 br_169 wl_81 vdd gnd cell_6t
Xbit_r82_c169 bl_169 br_169 wl_82 vdd gnd cell_6t
Xbit_r83_c169 bl_169 br_169 wl_83 vdd gnd cell_6t
Xbit_r84_c169 bl_169 br_169 wl_84 vdd gnd cell_6t
Xbit_r85_c169 bl_169 br_169 wl_85 vdd gnd cell_6t
Xbit_r86_c169 bl_169 br_169 wl_86 vdd gnd cell_6t
Xbit_r87_c169 bl_169 br_169 wl_87 vdd gnd cell_6t
Xbit_r88_c169 bl_169 br_169 wl_88 vdd gnd cell_6t
Xbit_r89_c169 bl_169 br_169 wl_89 vdd gnd cell_6t
Xbit_r90_c169 bl_169 br_169 wl_90 vdd gnd cell_6t
Xbit_r91_c169 bl_169 br_169 wl_91 vdd gnd cell_6t
Xbit_r92_c169 bl_169 br_169 wl_92 vdd gnd cell_6t
Xbit_r93_c169 bl_169 br_169 wl_93 vdd gnd cell_6t
Xbit_r94_c169 bl_169 br_169 wl_94 vdd gnd cell_6t
Xbit_r95_c169 bl_169 br_169 wl_95 vdd gnd cell_6t
Xbit_r96_c169 bl_169 br_169 wl_96 vdd gnd cell_6t
Xbit_r97_c169 bl_169 br_169 wl_97 vdd gnd cell_6t
Xbit_r98_c169 bl_169 br_169 wl_98 vdd gnd cell_6t
Xbit_r99_c169 bl_169 br_169 wl_99 vdd gnd cell_6t
Xbit_r100_c169 bl_169 br_169 wl_100 vdd gnd cell_6t
Xbit_r101_c169 bl_169 br_169 wl_101 vdd gnd cell_6t
Xbit_r102_c169 bl_169 br_169 wl_102 vdd gnd cell_6t
Xbit_r103_c169 bl_169 br_169 wl_103 vdd gnd cell_6t
Xbit_r104_c169 bl_169 br_169 wl_104 vdd gnd cell_6t
Xbit_r105_c169 bl_169 br_169 wl_105 vdd gnd cell_6t
Xbit_r106_c169 bl_169 br_169 wl_106 vdd gnd cell_6t
Xbit_r107_c169 bl_169 br_169 wl_107 vdd gnd cell_6t
Xbit_r108_c169 bl_169 br_169 wl_108 vdd gnd cell_6t
Xbit_r109_c169 bl_169 br_169 wl_109 vdd gnd cell_6t
Xbit_r110_c169 bl_169 br_169 wl_110 vdd gnd cell_6t
Xbit_r111_c169 bl_169 br_169 wl_111 vdd gnd cell_6t
Xbit_r112_c169 bl_169 br_169 wl_112 vdd gnd cell_6t
Xbit_r113_c169 bl_169 br_169 wl_113 vdd gnd cell_6t
Xbit_r114_c169 bl_169 br_169 wl_114 vdd gnd cell_6t
Xbit_r115_c169 bl_169 br_169 wl_115 vdd gnd cell_6t
Xbit_r116_c169 bl_169 br_169 wl_116 vdd gnd cell_6t
Xbit_r117_c169 bl_169 br_169 wl_117 vdd gnd cell_6t
Xbit_r118_c169 bl_169 br_169 wl_118 vdd gnd cell_6t
Xbit_r119_c169 bl_169 br_169 wl_119 vdd gnd cell_6t
Xbit_r120_c169 bl_169 br_169 wl_120 vdd gnd cell_6t
Xbit_r121_c169 bl_169 br_169 wl_121 vdd gnd cell_6t
Xbit_r122_c169 bl_169 br_169 wl_122 vdd gnd cell_6t
Xbit_r123_c169 bl_169 br_169 wl_123 vdd gnd cell_6t
Xbit_r124_c169 bl_169 br_169 wl_124 vdd gnd cell_6t
Xbit_r125_c169 bl_169 br_169 wl_125 vdd gnd cell_6t
Xbit_r126_c169 bl_169 br_169 wl_126 vdd gnd cell_6t
Xbit_r127_c169 bl_169 br_169 wl_127 vdd gnd cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd cell_6t
Xbit_r1_c170 bl_170 br_170 wl_1 vdd gnd cell_6t
Xbit_r2_c170 bl_170 br_170 wl_2 vdd gnd cell_6t
Xbit_r3_c170 bl_170 br_170 wl_3 vdd gnd cell_6t
Xbit_r4_c170 bl_170 br_170 wl_4 vdd gnd cell_6t
Xbit_r5_c170 bl_170 br_170 wl_5 vdd gnd cell_6t
Xbit_r6_c170 bl_170 br_170 wl_6 vdd gnd cell_6t
Xbit_r7_c170 bl_170 br_170 wl_7 vdd gnd cell_6t
Xbit_r8_c170 bl_170 br_170 wl_8 vdd gnd cell_6t
Xbit_r9_c170 bl_170 br_170 wl_9 vdd gnd cell_6t
Xbit_r10_c170 bl_170 br_170 wl_10 vdd gnd cell_6t
Xbit_r11_c170 bl_170 br_170 wl_11 vdd gnd cell_6t
Xbit_r12_c170 bl_170 br_170 wl_12 vdd gnd cell_6t
Xbit_r13_c170 bl_170 br_170 wl_13 vdd gnd cell_6t
Xbit_r14_c170 bl_170 br_170 wl_14 vdd gnd cell_6t
Xbit_r15_c170 bl_170 br_170 wl_15 vdd gnd cell_6t
Xbit_r16_c170 bl_170 br_170 wl_16 vdd gnd cell_6t
Xbit_r17_c170 bl_170 br_170 wl_17 vdd gnd cell_6t
Xbit_r18_c170 bl_170 br_170 wl_18 vdd gnd cell_6t
Xbit_r19_c170 bl_170 br_170 wl_19 vdd gnd cell_6t
Xbit_r20_c170 bl_170 br_170 wl_20 vdd gnd cell_6t
Xbit_r21_c170 bl_170 br_170 wl_21 vdd gnd cell_6t
Xbit_r22_c170 bl_170 br_170 wl_22 vdd gnd cell_6t
Xbit_r23_c170 bl_170 br_170 wl_23 vdd gnd cell_6t
Xbit_r24_c170 bl_170 br_170 wl_24 vdd gnd cell_6t
Xbit_r25_c170 bl_170 br_170 wl_25 vdd gnd cell_6t
Xbit_r26_c170 bl_170 br_170 wl_26 vdd gnd cell_6t
Xbit_r27_c170 bl_170 br_170 wl_27 vdd gnd cell_6t
Xbit_r28_c170 bl_170 br_170 wl_28 vdd gnd cell_6t
Xbit_r29_c170 bl_170 br_170 wl_29 vdd gnd cell_6t
Xbit_r30_c170 bl_170 br_170 wl_30 vdd gnd cell_6t
Xbit_r31_c170 bl_170 br_170 wl_31 vdd gnd cell_6t
Xbit_r32_c170 bl_170 br_170 wl_32 vdd gnd cell_6t
Xbit_r33_c170 bl_170 br_170 wl_33 vdd gnd cell_6t
Xbit_r34_c170 bl_170 br_170 wl_34 vdd gnd cell_6t
Xbit_r35_c170 bl_170 br_170 wl_35 vdd gnd cell_6t
Xbit_r36_c170 bl_170 br_170 wl_36 vdd gnd cell_6t
Xbit_r37_c170 bl_170 br_170 wl_37 vdd gnd cell_6t
Xbit_r38_c170 bl_170 br_170 wl_38 vdd gnd cell_6t
Xbit_r39_c170 bl_170 br_170 wl_39 vdd gnd cell_6t
Xbit_r40_c170 bl_170 br_170 wl_40 vdd gnd cell_6t
Xbit_r41_c170 bl_170 br_170 wl_41 vdd gnd cell_6t
Xbit_r42_c170 bl_170 br_170 wl_42 vdd gnd cell_6t
Xbit_r43_c170 bl_170 br_170 wl_43 vdd gnd cell_6t
Xbit_r44_c170 bl_170 br_170 wl_44 vdd gnd cell_6t
Xbit_r45_c170 bl_170 br_170 wl_45 vdd gnd cell_6t
Xbit_r46_c170 bl_170 br_170 wl_46 vdd gnd cell_6t
Xbit_r47_c170 bl_170 br_170 wl_47 vdd gnd cell_6t
Xbit_r48_c170 bl_170 br_170 wl_48 vdd gnd cell_6t
Xbit_r49_c170 bl_170 br_170 wl_49 vdd gnd cell_6t
Xbit_r50_c170 bl_170 br_170 wl_50 vdd gnd cell_6t
Xbit_r51_c170 bl_170 br_170 wl_51 vdd gnd cell_6t
Xbit_r52_c170 bl_170 br_170 wl_52 vdd gnd cell_6t
Xbit_r53_c170 bl_170 br_170 wl_53 vdd gnd cell_6t
Xbit_r54_c170 bl_170 br_170 wl_54 vdd gnd cell_6t
Xbit_r55_c170 bl_170 br_170 wl_55 vdd gnd cell_6t
Xbit_r56_c170 bl_170 br_170 wl_56 vdd gnd cell_6t
Xbit_r57_c170 bl_170 br_170 wl_57 vdd gnd cell_6t
Xbit_r58_c170 bl_170 br_170 wl_58 vdd gnd cell_6t
Xbit_r59_c170 bl_170 br_170 wl_59 vdd gnd cell_6t
Xbit_r60_c170 bl_170 br_170 wl_60 vdd gnd cell_6t
Xbit_r61_c170 bl_170 br_170 wl_61 vdd gnd cell_6t
Xbit_r62_c170 bl_170 br_170 wl_62 vdd gnd cell_6t
Xbit_r63_c170 bl_170 br_170 wl_63 vdd gnd cell_6t
Xbit_r64_c170 bl_170 br_170 wl_64 vdd gnd cell_6t
Xbit_r65_c170 bl_170 br_170 wl_65 vdd gnd cell_6t
Xbit_r66_c170 bl_170 br_170 wl_66 vdd gnd cell_6t
Xbit_r67_c170 bl_170 br_170 wl_67 vdd gnd cell_6t
Xbit_r68_c170 bl_170 br_170 wl_68 vdd gnd cell_6t
Xbit_r69_c170 bl_170 br_170 wl_69 vdd gnd cell_6t
Xbit_r70_c170 bl_170 br_170 wl_70 vdd gnd cell_6t
Xbit_r71_c170 bl_170 br_170 wl_71 vdd gnd cell_6t
Xbit_r72_c170 bl_170 br_170 wl_72 vdd gnd cell_6t
Xbit_r73_c170 bl_170 br_170 wl_73 vdd gnd cell_6t
Xbit_r74_c170 bl_170 br_170 wl_74 vdd gnd cell_6t
Xbit_r75_c170 bl_170 br_170 wl_75 vdd gnd cell_6t
Xbit_r76_c170 bl_170 br_170 wl_76 vdd gnd cell_6t
Xbit_r77_c170 bl_170 br_170 wl_77 vdd gnd cell_6t
Xbit_r78_c170 bl_170 br_170 wl_78 vdd gnd cell_6t
Xbit_r79_c170 bl_170 br_170 wl_79 vdd gnd cell_6t
Xbit_r80_c170 bl_170 br_170 wl_80 vdd gnd cell_6t
Xbit_r81_c170 bl_170 br_170 wl_81 vdd gnd cell_6t
Xbit_r82_c170 bl_170 br_170 wl_82 vdd gnd cell_6t
Xbit_r83_c170 bl_170 br_170 wl_83 vdd gnd cell_6t
Xbit_r84_c170 bl_170 br_170 wl_84 vdd gnd cell_6t
Xbit_r85_c170 bl_170 br_170 wl_85 vdd gnd cell_6t
Xbit_r86_c170 bl_170 br_170 wl_86 vdd gnd cell_6t
Xbit_r87_c170 bl_170 br_170 wl_87 vdd gnd cell_6t
Xbit_r88_c170 bl_170 br_170 wl_88 vdd gnd cell_6t
Xbit_r89_c170 bl_170 br_170 wl_89 vdd gnd cell_6t
Xbit_r90_c170 bl_170 br_170 wl_90 vdd gnd cell_6t
Xbit_r91_c170 bl_170 br_170 wl_91 vdd gnd cell_6t
Xbit_r92_c170 bl_170 br_170 wl_92 vdd gnd cell_6t
Xbit_r93_c170 bl_170 br_170 wl_93 vdd gnd cell_6t
Xbit_r94_c170 bl_170 br_170 wl_94 vdd gnd cell_6t
Xbit_r95_c170 bl_170 br_170 wl_95 vdd gnd cell_6t
Xbit_r96_c170 bl_170 br_170 wl_96 vdd gnd cell_6t
Xbit_r97_c170 bl_170 br_170 wl_97 vdd gnd cell_6t
Xbit_r98_c170 bl_170 br_170 wl_98 vdd gnd cell_6t
Xbit_r99_c170 bl_170 br_170 wl_99 vdd gnd cell_6t
Xbit_r100_c170 bl_170 br_170 wl_100 vdd gnd cell_6t
Xbit_r101_c170 bl_170 br_170 wl_101 vdd gnd cell_6t
Xbit_r102_c170 bl_170 br_170 wl_102 vdd gnd cell_6t
Xbit_r103_c170 bl_170 br_170 wl_103 vdd gnd cell_6t
Xbit_r104_c170 bl_170 br_170 wl_104 vdd gnd cell_6t
Xbit_r105_c170 bl_170 br_170 wl_105 vdd gnd cell_6t
Xbit_r106_c170 bl_170 br_170 wl_106 vdd gnd cell_6t
Xbit_r107_c170 bl_170 br_170 wl_107 vdd gnd cell_6t
Xbit_r108_c170 bl_170 br_170 wl_108 vdd gnd cell_6t
Xbit_r109_c170 bl_170 br_170 wl_109 vdd gnd cell_6t
Xbit_r110_c170 bl_170 br_170 wl_110 vdd gnd cell_6t
Xbit_r111_c170 bl_170 br_170 wl_111 vdd gnd cell_6t
Xbit_r112_c170 bl_170 br_170 wl_112 vdd gnd cell_6t
Xbit_r113_c170 bl_170 br_170 wl_113 vdd gnd cell_6t
Xbit_r114_c170 bl_170 br_170 wl_114 vdd gnd cell_6t
Xbit_r115_c170 bl_170 br_170 wl_115 vdd gnd cell_6t
Xbit_r116_c170 bl_170 br_170 wl_116 vdd gnd cell_6t
Xbit_r117_c170 bl_170 br_170 wl_117 vdd gnd cell_6t
Xbit_r118_c170 bl_170 br_170 wl_118 vdd gnd cell_6t
Xbit_r119_c170 bl_170 br_170 wl_119 vdd gnd cell_6t
Xbit_r120_c170 bl_170 br_170 wl_120 vdd gnd cell_6t
Xbit_r121_c170 bl_170 br_170 wl_121 vdd gnd cell_6t
Xbit_r122_c170 bl_170 br_170 wl_122 vdd gnd cell_6t
Xbit_r123_c170 bl_170 br_170 wl_123 vdd gnd cell_6t
Xbit_r124_c170 bl_170 br_170 wl_124 vdd gnd cell_6t
Xbit_r125_c170 bl_170 br_170 wl_125 vdd gnd cell_6t
Xbit_r126_c170 bl_170 br_170 wl_126 vdd gnd cell_6t
Xbit_r127_c170 bl_170 br_170 wl_127 vdd gnd cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd cell_6t
Xbit_r1_c171 bl_171 br_171 wl_1 vdd gnd cell_6t
Xbit_r2_c171 bl_171 br_171 wl_2 vdd gnd cell_6t
Xbit_r3_c171 bl_171 br_171 wl_3 vdd gnd cell_6t
Xbit_r4_c171 bl_171 br_171 wl_4 vdd gnd cell_6t
Xbit_r5_c171 bl_171 br_171 wl_5 vdd gnd cell_6t
Xbit_r6_c171 bl_171 br_171 wl_6 vdd gnd cell_6t
Xbit_r7_c171 bl_171 br_171 wl_7 vdd gnd cell_6t
Xbit_r8_c171 bl_171 br_171 wl_8 vdd gnd cell_6t
Xbit_r9_c171 bl_171 br_171 wl_9 vdd gnd cell_6t
Xbit_r10_c171 bl_171 br_171 wl_10 vdd gnd cell_6t
Xbit_r11_c171 bl_171 br_171 wl_11 vdd gnd cell_6t
Xbit_r12_c171 bl_171 br_171 wl_12 vdd gnd cell_6t
Xbit_r13_c171 bl_171 br_171 wl_13 vdd gnd cell_6t
Xbit_r14_c171 bl_171 br_171 wl_14 vdd gnd cell_6t
Xbit_r15_c171 bl_171 br_171 wl_15 vdd gnd cell_6t
Xbit_r16_c171 bl_171 br_171 wl_16 vdd gnd cell_6t
Xbit_r17_c171 bl_171 br_171 wl_17 vdd gnd cell_6t
Xbit_r18_c171 bl_171 br_171 wl_18 vdd gnd cell_6t
Xbit_r19_c171 bl_171 br_171 wl_19 vdd gnd cell_6t
Xbit_r20_c171 bl_171 br_171 wl_20 vdd gnd cell_6t
Xbit_r21_c171 bl_171 br_171 wl_21 vdd gnd cell_6t
Xbit_r22_c171 bl_171 br_171 wl_22 vdd gnd cell_6t
Xbit_r23_c171 bl_171 br_171 wl_23 vdd gnd cell_6t
Xbit_r24_c171 bl_171 br_171 wl_24 vdd gnd cell_6t
Xbit_r25_c171 bl_171 br_171 wl_25 vdd gnd cell_6t
Xbit_r26_c171 bl_171 br_171 wl_26 vdd gnd cell_6t
Xbit_r27_c171 bl_171 br_171 wl_27 vdd gnd cell_6t
Xbit_r28_c171 bl_171 br_171 wl_28 vdd gnd cell_6t
Xbit_r29_c171 bl_171 br_171 wl_29 vdd gnd cell_6t
Xbit_r30_c171 bl_171 br_171 wl_30 vdd gnd cell_6t
Xbit_r31_c171 bl_171 br_171 wl_31 vdd gnd cell_6t
Xbit_r32_c171 bl_171 br_171 wl_32 vdd gnd cell_6t
Xbit_r33_c171 bl_171 br_171 wl_33 vdd gnd cell_6t
Xbit_r34_c171 bl_171 br_171 wl_34 vdd gnd cell_6t
Xbit_r35_c171 bl_171 br_171 wl_35 vdd gnd cell_6t
Xbit_r36_c171 bl_171 br_171 wl_36 vdd gnd cell_6t
Xbit_r37_c171 bl_171 br_171 wl_37 vdd gnd cell_6t
Xbit_r38_c171 bl_171 br_171 wl_38 vdd gnd cell_6t
Xbit_r39_c171 bl_171 br_171 wl_39 vdd gnd cell_6t
Xbit_r40_c171 bl_171 br_171 wl_40 vdd gnd cell_6t
Xbit_r41_c171 bl_171 br_171 wl_41 vdd gnd cell_6t
Xbit_r42_c171 bl_171 br_171 wl_42 vdd gnd cell_6t
Xbit_r43_c171 bl_171 br_171 wl_43 vdd gnd cell_6t
Xbit_r44_c171 bl_171 br_171 wl_44 vdd gnd cell_6t
Xbit_r45_c171 bl_171 br_171 wl_45 vdd gnd cell_6t
Xbit_r46_c171 bl_171 br_171 wl_46 vdd gnd cell_6t
Xbit_r47_c171 bl_171 br_171 wl_47 vdd gnd cell_6t
Xbit_r48_c171 bl_171 br_171 wl_48 vdd gnd cell_6t
Xbit_r49_c171 bl_171 br_171 wl_49 vdd gnd cell_6t
Xbit_r50_c171 bl_171 br_171 wl_50 vdd gnd cell_6t
Xbit_r51_c171 bl_171 br_171 wl_51 vdd gnd cell_6t
Xbit_r52_c171 bl_171 br_171 wl_52 vdd gnd cell_6t
Xbit_r53_c171 bl_171 br_171 wl_53 vdd gnd cell_6t
Xbit_r54_c171 bl_171 br_171 wl_54 vdd gnd cell_6t
Xbit_r55_c171 bl_171 br_171 wl_55 vdd gnd cell_6t
Xbit_r56_c171 bl_171 br_171 wl_56 vdd gnd cell_6t
Xbit_r57_c171 bl_171 br_171 wl_57 vdd gnd cell_6t
Xbit_r58_c171 bl_171 br_171 wl_58 vdd gnd cell_6t
Xbit_r59_c171 bl_171 br_171 wl_59 vdd gnd cell_6t
Xbit_r60_c171 bl_171 br_171 wl_60 vdd gnd cell_6t
Xbit_r61_c171 bl_171 br_171 wl_61 vdd gnd cell_6t
Xbit_r62_c171 bl_171 br_171 wl_62 vdd gnd cell_6t
Xbit_r63_c171 bl_171 br_171 wl_63 vdd gnd cell_6t
Xbit_r64_c171 bl_171 br_171 wl_64 vdd gnd cell_6t
Xbit_r65_c171 bl_171 br_171 wl_65 vdd gnd cell_6t
Xbit_r66_c171 bl_171 br_171 wl_66 vdd gnd cell_6t
Xbit_r67_c171 bl_171 br_171 wl_67 vdd gnd cell_6t
Xbit_r68_c171 bl_171 br_171 wl_68 vdd gnd cell_6t
Xbit_r69_c171 bl_171 br_171 wl_69 vdd gnd cell_6t
Xbit_r70_c171 bl_171 br_171 wl_70 vdd gnd cell_6t
Xbit_r71_c171 bl_171 br_171 wl_71 vdd gnd cell_6t
Xbit_r72_c171 bl_171 br_171 wl_72 vdd gnd cell_6t
Xbit_r73_c171 bl_171 br_171 wl_73 vdd gnd cell_6t
Xbit_r74_c171 bl_171 br_171 wl_74 vdd gnd cell_6t
Xbit_r75_c171 bl_171 br_171 wl_75 vdd gnd cell_6t
Xbit_r76_c171 bl_171 br_171 wl_76 vdd gnd cell_6t
Xbit_r77_c171 bl_171 br_171 wl_77 vdd gnd cell_6t
Xbit_r78_c171 bl_171 br_171 wl_78 vdd gnd cell_6t
Xbit_r79_c171 bl_171 br_171 wl_79 vdd gnd cell_6t
Xbit_r80_c171 bl_171 br_171 wl_80 vdd gnd cell_6t
Xbit_r81_c171 bl_171 br_171 wl_81 vdd gnd cell_6t
Xbit_r82_c171 bl_171 br_171 wl_82 vdd gnd cell_6t
Xbit_r83_c171 bl_171 br_171 wl_83 vdd gnd cell_6t
Xbit_r84_c171 bl_171 br_171 wl_84 vdd gnd cell_6t
Xbit_r85_c171 bl_171 br_171 wl_85 vdd gnd cell_6t
Xbit_r86_c171 bl_171 br_171 wl_86 vdd gnd cell_6t
Xbit_r87_c171 bl_171 br_171 wl_87 vdd gnd cell_6t
Xbit_r88_c171 bl_171 br_171 wl_88 vdd gnd cell_6t
Xbit_r89_c171 bl_171 br_171 wl_89 vdd gnd cell_6t
Xbit_r90_c171 bl_171 br_171 wl_90 vdd gnd cell_6t
Xbit_r91_c171 bl_171 br_171 wl_91 vdd gnd cell_6t
Xbit_r92_c171 bl_171 br_171 wl_92 vdd gnd cell_6t
Xbit_r93_c171 bl_171 br_171 wl_93 vdd gnd cell_6t
Xbit_r94_c171 bl_171 br_171 wl_94 vdd gnd cell_6t
Xbit_r95_c171 bl_171 br_171 wl_95 vdd gnd cell_6t
Xbit_r96_c171 bl_171 br_171 wl_96 vdd gnd cell_6t
Xbit_r97_c171 bl_171 br_171 wl_97 vdd gnd cell_6t
Xbit_r98_c171 bl_171 br_171 wl_98 vdd gnd cell_6t
Xbit_r99_c171 bl_171 br_171 wl_99 vdd gnd cell_6t
Xbit_r100_c171 bl_171 br_171 wl_100 vdd gnd cell_6t
Xbit_r101_c171 bl_171 br_171 wl_101 vdd gnd cell_6t
Xbit_r102_c171 bl_171 br_171 wl_102 vdd gnd cell_6t
Xbit_r103_c171 bl_171 br_171 wl_103 vdd gnd cell_6t
Xbit_r104_c171 bl_171 br_171 wl_104 vdd gnd cell_6t
Xbit_r105_c171 bl_171 br_171 wl_105 vdd gnd cell_6t
Xbit_r106_c171 bl_171 br_171 wl_106 vdd gnd cell_6t
Xbit_r107_c171 bl_171 br_171 wl_107 vdd gnd cell_6t
Xbit_r108_c171 bl_171 br_171 wl_108 vdd gnd cell_6t
Xbit_r109_c171 bl_171 br_171 wl_109 vdd gnd cell_6t
Xbit_r110_c171 bl_171 br_171 wl_110 vdd gnd cell_6t
Xbit_r111_c171 bl_171 br_171 wl_111 vdd gnd cell_6t
Xbit_r112_c171 bl_171 br_171 wl_112 vdd gnd cell_6t
Xbit_r113_c171 bl_171 br_171 wl_113 vdd gnd cell_6t
Xbit_r114_c171 bl_171 br_171 wl_114 vdd gnd cell_6t
Xbit_r115_c171 bl_171 br_171 wl_115 vdd gnd cell_6t
Xbit_r116_c171 bl_171 br_171 wl_116 vdd gnd cell_6t
Xbit_r117_c171 bl_171 br_171 wl_117 vdd gnd cell_6t
Xbit_r118_c171 bl_171 br_171 wl_118 vdd gnd cell_6t
Xbit_r119_c171 bl_171 br_171 wl_119 vdd gnd cell_6t
Xbit_r120_c171 bl_171 br_171 wl_120 vdd gnd cell_6t
Xbit_r121_c171 bl_171 br_171 wl_121 vdd gnd cell_6t
Xbit_r122_c171 bl_171 br_171 wl_122 vdd gnd cell_6t
Xbit_r123_c171 bl_171 br_171 wl_123 vdd gnd cell_6t
Xbit_r124_c171 bl_171 br_171 wl_124 vdd gnd cell_6t
Xbit_r125_c171 bl_171 br_171 wl_125 vdd gnd cell_6t
Xbit_r126_c171 bl_171 br_171 wl_126 vdd gnd cell_6t
Xbit_r127_c171 bl_171 br_171 wl_127 vdd gnd cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd cell_6t
Xbit_r1_c172 bl_172 br_172 wl_1 vdd gnd cell_6t
Xbit_r2_c172 bl_172 br_172 wl_2 vdd gnd cell_6t
Xbit_r3_c172 bl_172 br_172 wl_3 vdd gnd cell_6t
Xbit_r4_c172 bl_172 br_172 wl_4 vdd gnd cell_6t
Xbit_r5_c172 bl_172 br_172 wl_5 vdd gnd cell_6t
Xbit_r6_c172 bl_172 br_172 wl_6 vdd gnd cell_6t
Xbit_r7_c172 bl_172 br_172 wl_7 vdd gnd cell_6t
Xbit_r8_c172 bl_172 br_172 wl_8 vdd gnd cell_6t
Xbit_r9_c172 bl_172 br_172 wl_9 vdd gnd cell_6t
Xbit_r10_c172 bl_172 br_172 wl_10 vdd gnd cell_6t
Xbit_r11_c172 bl_172 br_172 wl_11 vdd gnd cell_6t
Xbit_r12_c172 bl_172 br_172 wl_12 vdd gnd cell_6t
Xbit_r13_c172 bl_172 br_172 wl_13 vdd gnd cell_6t
Xbit_r14_c172 bl_172 br_172 wl_14 vdd gnd cell_6t
Xbit_r15_c172 bl_172 br_172 wl_15 vdd gnd cell_6t
Xbit_r16_c172 bl_172 br_172 wl_16 vdd gnd cell_6t
Xbit_r17_c172 bl_172 br_172 wl_17 vdd gnd cell_6t
Xbit_r18_c172 bl_172 br_172 wl_18 vdd gnd cell_6t
Xbit_r19_c172 bl_172 br_172 wl_19 vdd gnd cell_6t
Xbit_r20_c172 bl_172 br_172 wl_20 vdd gnd cell_6t
Xbit_r21_c172 bl_172 br_172 wl_21 vdd gnd cell_6t
Xbit_r22_c172 bl_172 br_172 wl_22 vdd gnd cell_6t
Xbit_r23_c172 bl_172 br_172 wl_23 vdd gnd cell_6t
Xbit_r24_c172 bl_172 br_172 wl_24 vdd gnd cell_6t
Xbit_r25_c172 bl_172 br_172 wl_25 vdd gnd cell_6t
Xbit_r26_c172 bl_172 br_172 wl_26 vdd gnd cell_6t
Xbit_r27_c172 bl_172 br_172 wl_27 vdd gnd cell_6t
Xbit_r28_c172 bl_172 br_172 wl_28 vdd gnd cell_6t
Xbit_r29_c172 bl_172 br_172 wl_29 vdd gnd cell_6t
Xbit_r30_c172 bl_172 br_172 wl_30 vdd gnd cell_6t
Xbit_r31_c172 bl_172 br_172 wl_31 vdd gnd cell_6t
Xbit_r32_c172 bl_172 br_172 wl_32 vdd gnd cell_6t
Xbit_r33_c172 bl_172 br_172 wl_33 vdd gnd cell_6t
Xbit_r34_c172 bl_172 br_172 wl_34 vdd gnd cell_6t
Xbit_r35_c172 bl_172 br_172 wl_35 vdd gnd cell_6t
Xbit_r36_c172 bl_172 br_172 wl_36 vdd gnd cell_6t
Xbit_r37_c172 bl_172 br_172 wl_37 vdd gnd cell_6t
Xbit_r38_c172 bl_172 br_172 wl_38 vdd gnd cell_6t
Xbit_r39_c172 bl_172 br_172 wl_39 vdd gnd cell_6t
Xbit_r40_c172 bl_172 br_172 wl_40 vdd gnd cell_6t
Xbit_r41_c172 bl_172 br_172 wl_41 vdd gnd cell_6t
Xbit_r42_c172 bl_172 br_172 wl_42 vdd gnd cell_6t
Xbit_r43_c172 bl_172 br_172 wl_43 vdd gnd cell_6t
Xbit_r44_c172 bl_172 br_172 wl_44 vdd gnd cell_6t
Xbit_r45_c172 bl_172 br_172 wl_45 vdd gnd cell_6t
Xbit_r46_c172 bl_172 br_172 wl_46 vdd gnd cell_6t
Xbit_r47_c172 bl_172 br_172 wl_47 vdd gnd cell_6t
Xbit_r48_c172 bl_172 br_172 wl_48 vdd gnd cell_6t
Xbit_r49_c172 bl_172 br_172 wl_49 vdd gnd cell_6t
Xbit_r50_c172 bl_172 br_172 wl_50 vdd gnd cell_6t
Xbit_r51_c172 bl_172 br_172 wl_51 vdd gnd cell_6t
Xbit_r52_c172 bl_172 br_172 wl_52 vdd gnd cell_6t
Xbit_r53_c172 bl_172 br_172 wl_53 vdd gnd cell_6t
Xbit_r54_c172 bl_172 br_172 wl_54 vdd gnd cell_6t
Xbit_r55_c172 bl_172 br_172 wl_55 vdd gnd cell_6t
Xbit_r56_c172 bl_172 br_172 wl_56 vdd gnd cell_6t
Xbit_r57_c172 bl_172 br_172 wl_57 vdd gnd cell_6t
Xbit_r58_c172 bl_172 br_172 wl_58 vdd gnd cell_6t
Xbit_r59_c172 bl_172 br_172 wl_59 vdd gnd cell_6t
Xbit_r60_c172 bl_172 br_172 wl_60 vdd gnd cell_6t
Xbit_r61_c172 bl_172 br_172 wl_61 vdd gnd cell_6t
Xbit_r62_c172 bl_172 br_172 wl_62 vdd gnd cell_6t
Xbit_r63_c172 bl_172 br_172 wl_63 vdd gnd cell_6t
Xbit_r64_c172 bl_172 br_172 wl_64 vdd gnd cell_6t
Xbit_r65_c172 bl_172 br_172 wl_65 vdd gnd cell_6t
Xbit_r66_c172 bl_172 br_172 wl_66 vdd gnd cell_6t
Xbit_r67_c172 bl_172 br_172 wl_67 vdd gnd cell_6t
Xbit_r68_c172 bl_172 br_172 wl_68 vdd gnd cell_6t
Xbit_r69_c172 bl_172 br_172 wl_69 vdd gnd cell_6t
Xbit_r70_c172 bl_172 br_172 wl_70 vdd gnd cell_6t
Xbit_r71_c172 bl_172 br_172 wl_71 vdd gnd cell_6t
Xbit_r72_c172 bl_172 br_172 wl_72 vdd gnd cell_6t
Xbit_r73_c172 bl_172 br_172 wl_73 vdd gnd cell_6t
Xbit_r74_c172 bl_172 br_172 wl_74 vdd gnd cell_6t
Xbit_r75_c172 bl_172 br_172 wl_75 vdd gnd cell_6t
Xbit_r76_c172 bl_172 br_172 wl_76 vdd gnd cell_6t
Xbit_r77_c172 bl_172 br_172 wl_77 vdd gnd cell_6t
Xbit_r78_c172 bl_172 br_172 wl_78 vdd gnd cell_6t
Xbit_r79_c172 bl_172 br_172 wl_79 vdd gnd cell_6t
Xbit_r80_c172 bl_172 br_172 wl_80 vdd gnd cell_6t
Xbit_r81_c172 bl_172 br_172 wl_81 vdd gnd cell_6t
Xbit_r82_c172 bl_172 br_172 wl_82 vdd gnd cell_6t
Xbit_r83_c172 bl_172 br_172 wl_83 vdd gnd cell_6t
Xbit_r84_c172 bl_172 br_172 wl_84 vdd gnd cell_6t
Xbit_r85_c172 bl_172 br_172 wl_85 vdd gnd cell_6t
Xbit_r86_c172 bl_172 br_172 wl_86 vdd gnd cell_6t
Xbit_r87_c172 bl_172 br_172 wl_87 vdd gnd cell_6t
Xbit_r88_c172 bl_172 br_172 wl_88 vdd gnd cell_6t
Xbit_r89_c172 bl_172 br_172 wl_89 vdd gnd cell_6t
Xbit_r90_c172 bl_172 br_172 wl_90 vdd gnd cell_6t
Xbit_r91_c172 bl_172 br_172 wl_91 vdd gnd cell_6t
Xbit_r92_c172 bl_172 br_172 wl_92 vdd gnd cell_6t
Xbit_r93_c172 bl_172 br_172 wl_93 vdd gnd cell_6t
Xbit_r94_c172 bl_172 br_172 wl_94 vdd gnd cell_6t
Xbit_r95_c172 bl_172 br_172 wl_95 vdd gnd cell_6t
Xbit_r96_c172 bl_172 br_172 wl_96 vdd gnd cell_6t
Xbit_r97_c172 bl_172 br_172 wl_97 vdd gnd cell_6t
Xbit_r98_c172 bl_172 br_172 wl_98 vdd gnd cell_6t
Xbit_r99_c172 bl_172 br_172 wl_99 vdd gnd cell_6t
Xbit_r100_c172 bl_172 br_172 wl_100 vdd gnd cell_6t
Xbit_r101_c172 bl_172 br_172 wl_101 vdd gnd cell_6t
Xbit_r102_c172 bl_172 br_172 wl_102 vdd gnd cell_6t
Xbit_r103_c172 bl_172 br_172 wl_103 vdd gnd cell_6t
Xbit_r104_c172 bl_172 br_172 wl_104 vdd gnd cell_6t
Xbit_r105_c172 bl_172 br_172 wl_105 vdd gnd cell_6t
Xbit_r106_c172 bl_172 br_172 wl_106 vdd gnd cell_6t
Xbit_r107_c172 bl_172 br_172 wl_107 vdd gnd cell_6t
Xbit_r108_c172 bl_172 br_172 wl_108 vdd gnd cell_6t
Xbit_r109_c172 bl_172 br_172 wl_109 vdd gnd cell_6t
Xbit_r110_c172 bl_172 br_172 wl_110 vdd gnd cell_6t
Xbit_r111_c172 bl_172 br_172 wl_111 vdd gnd cell_6t
Xbit_r112_c172 bl_172 br_172 wl_112 vdd gnd cell_6t
Xbit_r113_c172 bl_172 br_172 wl_113 vdd gnd cell_6t
Xbit_r114_c172 bl_172 br_172 wl_114 vdd gnd cell_6t
Xbit_r115_c172 bl_172 br_172 wl_115 vdd gnd cell_6t
Xbit_r116_c172 bl_172 br_172 wl_116 vdd gnd cell_6t
Xbit_r117_c172 bl_172 br_172 wl_117 vdd gnd cell_6t
Xbit_r118_c172 bl_172 br_172 wl_118 vdd gnd cell_6t
Xbit_r119_c172 bl_172 br_172 wl_119 vdd gnd cell_6t
Xbit_r120_c172 bl_172 br_172 wl_120 vdd gnd cell_6t
Xbit_r121_c172 bl_172 br_172 wl_121 vdd gnd cell_6t
Xbit_r122_c172 bl_172 br_172 wl_122 vdd gnd cell_6t
Xbit_r123_c172 bl_172 br_172 wl_123 vdd gnd cell_6t
Xbit_r124_c172 bl_172 br_172 wl_124 vdd gnd cell_6t
Xbit_r125_c172 bl_172 br_172 wl_125 vdd gnd cell_6t
Xbit_r126_c172 bl_172 br_172 wl_126 vdd gnd cell_6t
Xbit_r127_c172 bl_172 br_172 wl_127 vdd gnd cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd cell_6t
Xbit_r1_c173 bl_173 br_173 wl_1 vdd gnd cell_6t
Xbit_r2_c173 bl_173 br_173 wl_2 vdd gnd cell_6t
Xbit_r3_c173 bl_173 br_173 wl_3 vdd gnd cell_6t
Xbit_r4_c173 bl_173 br_173 wl_4 vdd gnd cell_6t
Xbit_r5_c173 bl_173 br_173 wl_5 vdd gnd cell_6t
Xbit_r6_c173 bl_173 br_173 wl_6 vdd gnd cell_6t
Xbit_r7_c173 bl_173 br_173 wl_7 vdd gnd cell_6t
Xbit_r8_c173 bl_173 br_173 wl_8 vdd gnd cell_6t
Xbit_r9_c173 bl_173 br_173 wl_9 vdd gnd cell_6t
Xbit_r10_c173 bl_173 br_173 wl_10 vdd gnd cell_6t
Xbit_r11_c173 bl_173 br_173 wl_11 vdd gnd cell_6t
Xbit_r12_c173 bl_173 br_173 wl_12 vdd gnd cell_6t
Xbit_r13_c173 bl_173 br_173 wl_13 vdd gnd cell_6t
Xbit_r14_c173 bl_173 br_173 wl_14 vdd gnd cell_6t
Xbit_r15_c173 bl_173 br_173 wl_15 vdd gnd cell_6t
Xbit_r16_c173 bl_173 br_173 wl_16 vdd gnd cell_6t
Xbit_r17_c173 bl_173 br_173 wl_17 vdd gnd cell_6t
Xbit_r18_c173 bl_173 br_173 wl_18 vdd gnd cell_6t
Xbit_r19_c173 bl_173 br_173 wl_19 vdd gnd cell_6t
Xbit_r20_c173 bl_173 br_173 wl_20 vdd gnd cell_6t
Xbit_r21_c173 bl_173 br_173 wl_21 vdd gnd cell_6t
Xbit_r22_c173 bl_173 br_173 wl_22 vdd gnd cell_6t
Xbit_r23_c173 bl_173 br_173 wl_23 vdd gnd cell_6t
Xbit_r24_c173 bl_173 br_173 wl_24 vdd gnd cell_6t
Xbit_r25_c173 bl_173 br_173 wl_25 vdd gnd cell_6t
Xbit_r26_c173 bl_173 br_173 wl_26 vdd gnd cell_6t
Xbit_r27_c173 bl_173 br_173 wl_27 vdd gnd cell_6t
Xbit_r28_c173 bl_173 br_173 wl_28 vdd gnd cell_6t
Xbit_r29_c173 bl_173 br_173 wl_29 vdd gnd cell_6t
Xbit_r30_c173 bl_173 br_173 wl_30 vdd gnd cell_6t
Xbit_r31_c173 bl_173 br_173 wl_31 vdd gnd cell_6t
Xbit_r32_c173 bl_173 br_173 wl_32 vdd gnd cell_6t
Xbit_r33_c173 bl_173 br_173 wl_33 vdd gnd cell_6t
Xbit_r34_c173 bl_173 br_173 wl_34 vdd gnd cell_6t
Xbit_r35_c173 bl_173 br_173 wl_35 vdd gnd cell_6t
Xbit_r36_c173 bl_173 br_173 wl_36 vdd gnd cell_6t
Xbit_r37_c173 bl_173 br_173 wl_37 vdd gnd cell_6t
Xbit_r38_c173 bl_173 br_173 wl_38 vdd gnd cell_6t
Xbit_r39_c173 bl_173 br_173 wl_39 vdd gnd cell_6t
Xbit_r40_c173 bl_173 br_173 wl_40 vdd gnd cell_6t
Xbit_r41_c173 bl_173 br_173 wl_41 vdd gnd cell_6t
Xbit_r42_c173 bl_173 br_173 wl_42 vdd gnd cell_6t
Xbit_r43_c173 bl_173 br_173 wl_43 vdd gnd cell_6t
Xbit_r44_c173 bl_173 br_173 wl_44 vdd gnd cell_6t
Xbit_r45_c173 bl_173 br_173 wl_45 vdd gnd cell_6t
Xbit_r46_c173 bl_173 br_173 wl_46 vdd gnd cell_6t
Xbit_r47_c173 bl_173 br_173 wl_47 vdd gnd cell_6t
Xbit_r48_c173 bl_173 br_173 wl_48 vdd gnd cell_6t
Xbit_r49_c173 bl_173 br_173 wl_49 vdd gnd cell_6t
Xbit_r50_c173 bl_173 br_173 wl_50 vdd gnd cell_6t
Xbit_r51_c173 bl_173 br_173 wl_51 vdd gnd cell_6t
Xbit_r52_c173 bl_173 br_173 wl_52 vdd gnd cell_6t
Xbit_r53_c173 bl_173 br_173 wl_53 vdd gnd cell_6t
Xbit_r54_c173 bl_173 br_173 wl_54 vdd gnd cell_6t
Xbit_r55_c173 bl_173 br_173 wl_55 vdd gnd cell_6t
Xbit_r56_c173 bl_173 br_173 wl_56 vdd gnd cell_6t
Xbit_r57_c173 bl_173 br_173 wl_57 vdd gnd cell_6t
Xbit_r58_c173 bl_173 br_173 wl_58 vdd gnd cell_6t
Xbit_r59_c173 bl_173 br_173 wl_59 vdd gnd cell_6t
Xbit_r60_c173 bl_173 br_173 wl_60 vdd gnd cell_6t
Xbit_r61_c173 bl_173 br_173 wl_61 vdd gnd cell_6t
Xbit_r62_c173 bl_173 br_173 wl_62 vdd gnd cell_6t
Xbit_r63_c173 bl_173 br_173 wl_63 vdd gnd cell_6t
Xbit_r64_c173 bl_173 br_173 wl_64 vdd gnd cell_6t
Xbit_r65_c173 bl_173 br_173 wl_65 vdd gnd cell_6t
Xbit_r66_c173 bl_173 br_173 wl_66 vdd gnd cell_6t
Xbit_r67_c173 bl_173 br_173 wl_67 vdd gnd cell_6t
Xbit_r68_c173 bl_173 br_173 wl_68 vdd gnd cell_6t
Xbit_r69_c173 bl_173 br_173 wl_69 vdd gnd cell_6t
Xbit_r70_c173 bl_173 br_173 wl_70 vdd gnd cell_6t
Xbit_r71_c173 bl_173 br_173 wl_71 vdd gnd cell_6t
Xbit_r72_c173 bl_173 br_173 wl_72 vdd gnd cell_6t
Xbit_r73_c173 bl_173 br_173 wl_73 vdd gnd cell_6t
Xbit_r74_c173 bl_173 br_173 wl_74 vdd gnd cell_6t
Xbit_r75_c173 bl_173 br_173 wl_75 vdd gnd cell_6t
Xbit_r76_c173 bl_173 br_173 wl_76 vdd gnd cell_6t
Xbit_r77_c173 bl_173 br_173 wl_77 vdd gnd cell_6t
Xbit_r78_c173 bl_173 br_173 wl_78 vdd gnd cell_6t
Xbit_r79_c173 bl_173 br_173 wl_79 vdd gnd cell_6t
Xbit_r80_c173 bl_173 br_173 wl_80 vdd gnd cell_6t
Xbit_r81_c173 bl_173 br_173 wl_81 vdd gnd cell_6t
Xbit_r82_c173 bl_173 br_173 wl_82 vdd gnd cell_6t
Xbit_r83_c173 bl_173 br_173 wl_83 vdd gnd cell_6t
Xbit_r84_c173 bl_173 br_173 wl_84 vdd gnd cell_6t
Xbit_r85_c173 bl_173 br_173 wl_85 vdd gnd cell_6t
Xbit_r86_c173 bl_173 br_173 wl_86 vdd gnd cell_6t
Xbit_r87_c173 bl_173 br_173 wl_87 vdd gnd cell_6t
Xbit_r88_c173 bl_173 br_173 wl_88 vdd gnd cell_6t
Xbit_r89_c173 bl_173 br_173 wl_89 vdd gnd cell_6t
Xbit_r90_c173 bl_173 br_173 wl_90 vdd gnd cell_6t
Xbit_r91_c173 bl_173 br_173 wl_91 vdd gnd cell_6t
Xbit_r92_c173 bl_173 br_173 wl_92 vdd gnd cell_6t
Xbit_r93_c173 bl_173 br_173 wl_93 vdd gnd cell_6t
Xbit_r94_c173 bl_173 br_173 wl_94 vdd gnd cell_6t
Xbit_r95_c173 bl_173 br_173 wl_95 vdd gnd cell_6t
Xbit_r96_c173 bl_173 br_173 wl_96 vdd gnd cell_6t
Xbit_r97_c173 bl_173 br_173 wl_97 vdd gnd cell_6t
Xbit_r98_c173 bl_173 br_173 wl_98 vdd gnd cell_6t
Xbit_r99_c173 bl_173 br_173 wl_99 vdd gnd cell_6t
Xbit_r100_c173 bl_173 br_173 wl_100 vdd gnd cell_6t
Xbit_r101_c173 bl_173 br_173 wl_101 vdd gnd cell_6t
Xbit_r102_c173 bl_173 br_173 wl_102 vdd gnd cell_6t
Xbit_r103_c173 bl_173 br_173 wl_103 vdd gnd cell_6t
Xbit_r104_c173 bl_173 br_173 wl_104 vdd gnd cell_6t
Xbit_r105_c173 bl_173 br_173 wl_105 vdd gnd cell_6t
Xbit_r106_c173 bl_173 br_173 wl_106 vdd gnd cell_6t
Xbit_r107_c173 bl_173 br_173 wl_107 vdd gnd cell_6t
Xbit_r108_c173 bl_173 br_173 wl_108 vdd gnd cell_6t
Xbit_r109_c173 bl_173 br_173 wl_109 vdd gnd cell_6t
Xbit_r110_c173 bl_173 br_173 wl_110 vdd gnd cell_6t
Xbit_r111_c173 bl_173 br_173 wl_111 vdd gnd cell_6t
Xbit_r112_c173 bl_173 br_173 wl_112 vdd gnd cell_6t
Xbit_r113_c173 bl_173 br_173 wl_113 vdd gnd cell_6t
Xbit_r114_c173 bl_173 br_173 wl_114 vdd gnd cell_6t
Xbit_r115_c173 bl_173 br_173 wl_115 vdd gnd cell_6t
Xbit_r116_c173 bl_173 br_173 wl_116 vdd gnd cell_6t
Xbit_r117_c173 bl_173 br_173 wl_117 vdd gnd cell_6t
Xbit_r118_c173 bl_173 br_173 wl_118 vdd gnd cell_6t
Xbit_r119_c173 bl_173 br_173 wl_119 vdd gnd cell_6t
Xbit_r120_c173 bl_173 br_173 wl_120 vdd gnd cell_6t
Xbit_r121_c173 bl_173 br_173 wl_121 vdd gnd cell_6t
Xbit_r122_c173 bl_173 br_173 wl_122 vdd gnd cell_6t
Xbit_r123_c173 bl_173 br_173 wl_123 vdd gnd cell_6t
Xbit_r124_c173 bl_173 br_173 wl_124 vdd gnd cell_6t
Xbit_r125_c173 bl_173 br_173 wl_125 vdd gnd cell_6t
Xbit_r126_c173 bl_173 br_173 wl_126 vdd gnd cell_6t
Xbit_r127_c173 bl_173 br_173 wl_127 vdd gnd cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd cell_6t
Xbit_r1_c174 bl_174 br_174 wl_1 vdd gnd cell_6t
Xbit_r2_c174 bl_174 br_174 wl_2 vdd gnd cell_6t
Xbit_r3_c174 bl_174 br_174 wl_3 vdd gnd cell_6t
Xbit_r4_c174 bl_174 br_174 wl_4 vdd gnd cell_6t
Xbit_r5_c174 bl_174 br_174 wl_5 vdd gnd cell_6t
Xbit_r6_c174 bl_174 br_174 wl_6 vdd gnd cell_6t
Xbit_r7_c174 bl_174 br_174 wl_7 vdd gnd cell_6t
Xbit_r8_c174 bl_174 br_174 wl_8 vdd gnd cell_6t
Xbit_r9_c174 bl_174 br_174 wl_9 vdd gnd cell_6t
Xbit_r10_c174 bl_174 br_174 wl_10 vdd gnd cell_6t
Xbit_r11_c174 bl_174 br_174 wl_11 vdd gnd cell_6t
Xbit_r12_c174 bl_174 br_174 wl_12 vdd gnd cell_6t
Xbit_r13_c174 bl_174 br_174 wl_13 vdd gnd cell_6t
Xbit_r14_c174 bl_174 br_174 wl_14 vdd gnd cell_6t
Xbit_r15_c174 bl_174 br_174 wl_15 vdd gnd cell_6t
Xbit_r16_c174 bl_174 br_174 wl_16 vdd gnd cell_6t
Xbit_r17_c174 bl_174 br_174 wl_17 vdd gnd cell_6t
Xbit_r18_c174 bl_174 br_174 wl_18 vdd gnd cell_6t
Xbit_r19_c174 bl_174 br_174 wl_19 vdd gnd cell_6t
Xbit_r20_c174 bl_174 br_174 wl_20 vdd gnd cell_6t
Xbit_r21_c174 bl_174 br_174 wl_21 vdd gnd cell_6t
Xbit_r22_c174 bl_174 br_174 wl_22 vdd gnd cell_6t
Xbit_r23_c174 bl_174 br_174 wl_23 vdd gnd cell_6t
Xbit_r24_c174 bl_174 br_174 wl_24 vdd gnd cell_6t
Xbit_r25_c174 bl_174 br_174 wl_25 vdd gnd cell_6t
Xbit_r26_c174 bl_174 br_174 wl_26 vdd gnd cell_6t
Xbit_r27_c174 bl_174 br_174 wl_27 vdd gnd cell_6t
Xbit_r28_c174 bl_174 br_174 wl_28 vdd gnd cell_6t
Xbit_r29_c174 bl_174 br_174 wl_29 vdd gnd cell_6t
Xbit_r30_c174 bl_174 br_174 wl_30 vdd gnd cell_6t
Xbit_r31_c174 bl_174 br_174 wl_31 vdd gnd cell_6t
Xbit_r32_c174 bl_174 br_174 wl_32 vdd gnd cell_6t
Xbit_r33_c174 bl_174 br_174 wl_33 vdd gnd cell_6t
Xbit_r34_c174 bl_174 br_174 wl_34 vdd gnd cell_6t
Xbit_r35_c174 bl_174 br_174 wl_35 vdd gnd cell_6t
Xbit_r36_c174 bl_174 br_174 wl_36 vdd gnd cell_6t
Xbit_r37_c174 bl_174 br_174 wl_37 vdd gnd cell_6t
Xbit_r38_c174 bl_174 br_174 wl_38 vdd gnd cell_6t
Xbit_r39_c174 bl_174 br_174 wl_39 vdd gnd cell_6t
Xbit_r40_c174 bl_174 br_174 wl_40 vdd gnd cell_6t
Xbit_r41_c174 bl_174 br_174 wl_41 vdd gnd cell_6t
Xbit_r42_c174 bl_174 br_174 wl_42 vdd gnd cell_6t
Xbit_r43_c174 bl_174 br_174 wl_43 vdd gnd cell_6t
Xbit_r44_c174 bl_174 br_174 wl_44 vdd gnd cell_6t
Xbit_r45_c174 bl_174 br_174 wl_45 vdd gnd cell_6t
Xbit_r46_c174 bl_174 br_174 wl_46 vdd gnd cell_6t
Xbit_r47_c174 bl_174 br_174 wl_47 vdd gnd cell_6t
Xbit_r48_c174 bl_174 br_174 wl_48 vdd gnd cell_6t
Xbit_r49_c174 bl_174 br_174 wl_49 vdd gnd cell_6t
Xbit_r50_c174 bl_174 br_174 wl_50 vdd gnd cell_6t
Xbit_r51_c174 bl_174 br_174 wl_51 vdd gnd cell_6t
Xbit_r52_c174 bl_174 br_174 wl_52 vdd gnd cell_6t
Xbit_r53_c174 bl_174 br_174 wl_53 vdd gnd cell_6t
Xbit_r54_c174 bl_174 br_174 wl_54 vdd gnd cell_6t
Xbit_r55_c174 bl_174 br_174 wl_55 vdd gnd cell_6t
Xbit_r56_c174 bl_174 br_174 wl_56 vdd gnd cell_6t
Xbit_r57_c174 bl_174 br_174 wl_57 vdd gnd cell_6t
Xbit_r58_c174 bl_174 br_174 wl_58 vdd gnd cell_6t
Xbit_r59_c174 bl_174 br_174 wl_59 vdd gnd cell_6t
Xbit_r60_c174 bl_174 br_174 wl_60 vdd gnd cell_6t
Xbit_r61_c174 bl_174 br_174 wl_61 vdd gnd cell_6t
Xbit_r62_c174 bl_174 br_174 wl_62 vdd gnd cell_6t
Xbit_r63_c174 bl_174 br_174 wl_63 vdd gnd cell_6t
Xbit_r64_c174 bl_174 br_174 wl_64 vdd gnd cell_6t
Xbit_r65_c174 bl_174 br_174 wl_65 vdd gnd cell_6t
Xbit_r66_c174 bl_174 br_174 wl_66 vdd gnd cell_6t
Xbit_r67_c174 bl_174 br_174 wl_67 vdd gnd cell_6t
Xbit_r68_c174 bl_174 br_174 wl_68 vdd gnd cell_6t
Xbit_r69_c174 bl_174 br_174 wl_69 vdd gnd cell_6t
Xbit_r70_c174 bl_174 br_174 wl_70 vdd gnd cell_6t
Xbit_r71_c174 bl_174 br_174 wl_71 vdd gnd cell_6t
Xbit_r72_c174 bl_174 br_174 wl_72 vdd gnd cell_6t
Xbit_r73_c174 bl_174 br_174 wl_73 vdd gnd cell_6t
Xbit_r74_c174 bl_174 br_174 wl_74 vdd gnd cell_6t
Xbit_r75_c174 bl_174 br_174 wl_75 vdd gnd cell_6t
Xbit_r76_c174 bl_174 br_174 wl_76 vdd gnd cell_6t
Xbit_r77_c174 bl_174 br_174 wl_77 vdd gnd cell_6t
Xbit_r78_c174 bl_174 br_174 wl_78 vdd gnd cell_6t
Xbit_r79_c174 bl_174 br_174 wl_79 vdd gnd cell_6t
Xbit_r80_c174 bl_174 br_174 wl_80 vdd gnd cell_6t
Xbit_r81_c174 bl_174 br_174 wl_81 vdd gnd cell_6t
Xbit_r82_c174 bl_174 br_174 wl_82 vdd gnd cell_6t
Xbit_r83_c174 bl_174 br_174 wl_83 vdd gnd cell_6t
Xbit_r84_c174 bl_174 br_174 wl_84 vdd gnd cell_6t
Xbit_r85_c174 bl_174 br_174 wl_85 vdd gnd cell_6t
Xbit_r86_c174 bl_174 br_174 wl_86 vdd gnd cell_6t
Xbit_r87_c174 bl_174 br_174 wl_87 vdd gnd cell_6t
Xbit_r88_c174 bl_174 br_174 wl_88 vdd gnd cell_6t
Xbit_r89_c174 bl_174 br_174 wl_89 vdd gnd cell_6t
Xbit_r90_c174 bl_174 br_174 wl_90 vdd gnd cell_6t
Xbit_r91_c174 bl_174 br_174 wl_91 vdd gnd cell_6t
Xbit_r92_c174 bl_174 br_174 wl_92 vdd gnd cell_6t
Xbit_r93_c174 bl_174 br_174 wl_93 vdd gnd cell_6t
Xbit_r94_c174 bl_174 br_174 wl_94 vdd gnd cell_6t
Xbit_r95_c174 bl_174 br_174 wl_95 vdd gnd cell_6t
Xbit_r96_c174 bl_174 br_174 wl_96 vdd gnd cell_6t
Xbit_r97_c174 bl_174 br_174 wl_97 vdd gnd cell_6t
Xbit_r98_c174 bl_174 br_174 wl_98 vdd gnd cell_6t
Xbit_r99_c174 bl_174 br_174 wl_99 vdd gnd cell_6t
Xbit_r100_c174 bl_174 br_174 wl_100 vdd gnd cell_6t
Xbit_r101_c174 bl_174 br_174 wl_101 vdd gnd cell_6t
Xbit_r102_c174 bl_174 br_174 wl_102 vdd gnd cell_6t
Xbit_r103_c174 bl_174 br_174 wl_103 vdd gnd cell_6t
Xbit_r104_c174 bl_174 br_174 wl_104 vdd gnd cell_6t
Xbit_r105_c174 bl_174 br_174 wl_105 vdd gnd cell_6t
Xbit_r106_c174 bl_174 br_174 wl_106 vdd gnd cell_6t
Xbit_r107_c174 bl_174 br_174 wl_107 vdd gnd cell_6t
Xbit_r108_c174 bl_174 br_174 wl_108 vdd gnd cell_6t
Xbit_r109_c174 bl_174 br_174 wl_109 vdd gnd cell_6t
Xbit_r110_c174 bl_174 br_174 wl_110 vdd gnd cell_6t
Xbit_r111_c174 bl_174 br_174 wl_111 vdd gnd cell_6t
Xbit_r112_c174 bl_174 br_174 wl_112 vdd gnd cell_6t
Xbit_r113_c174 bl_174 br_174 wl_113 vdd gnd cell_6t
Xbit_r114_c174 bl_174 br_174 wl_114 vdd gnd cell_6t
Xbit_r115_c174 bl_174 br_174 wl_115 vdd gnd cell_6t
Xbit_r116_c174 bl_174 br_174 wl_116 vdd gnd cell_6t
Xbit_r117_c174 bl_174 br_174 wl_117 vdd gnd cell_6t
Xbit_r118_c174 bl_174 br_174 wl_118 vdd gnd cell_6t
Xbit_r119_c174 bl_174 br_174 wl_119 vdd gnd cell_6t
Xbit_r120_c174 bl_174 br_174 wl_120 vdd gnd cell_6t
Xbit_r121_c174 bl_174 br_174 wl_121 vdd gnd cell_6t
Xbit_r122_c174 bl_174 br_174 wl_122 vdd gnd cell_6t
Xbit_r123_c174 bl_174 br_174 wl_123 vdd gnd cell_6t
Xbit_r124_c174 bl_174 br_174 wl_124 vdd gnd cell_6t
Xbit_r125_c174 bl_174 br_174 wl_125 vdd gnd cell_6t
Xbit_r126_c174 bl_174 br_174 wl_126 vdd gnd cell_6t
Xbit_r127_c174 bl_174 br_174 wl_127 vdd gnd cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd cell_6t
Xbit_r1_c175 bl_175 br_175 wl_1 vdd gnd cell_6t
Xbit_r2_c175 bl_175 br_175 wl_2 vdd gnd cell_6t
Xbit_r3_c175 bl_175 br_175 wl_3 vdd gnd cell_6t
Xbit_r4_c175 bl_175 br_175 wl_4 vdd gnd cell_6t
Xbit_r5_c175 bl_175 br_175 wl_5 vdd gnd cell_6t
Xbit_r6_c175 bl_175 br_175 wl_6 vdd gnd cell_6t
Xbit_r7_c175 bl_175 br_175 wl_7 vdd gnd cell_6t
Xbit_r8_c175 bl_175 br_175 wl_8 vdd gnd cell_6t
Xbit_r9_c175 bl_175 br_175 wl_9 vdd gnd cell_6t
Xbit_r10_c175 bl_175 br_175 wl_10 vdd gnd cell_6t
Xbit_r11_c175 bl_175 br_175 wl_11 vdd gnd cell_6t
Xbit_r12_c175 bl_175 br_175 wl_12 vdd gnd cell_6t
Xbit_r13_c175 bl_175 br_175 wl_13 vdd gnd cell_6t
Xbit_r14_c175 bl_175 br_175 wl_14 vdd gnd cell_6t
Xbit_r15_c175 bl_175 br_175 wl_15 vdd gnd cell_6t
Xbit_r16_c175 bl_175 br_175 wl_16 vdd gnd cell_6t
Xbit_r17_c175 bl_175 br_175 wl_17 vdd gnd cell_6t
Xbit_r18_c175 bl_175 br_175 wl_18 vdd gnd cell_6t
Xbit_r19_c175 bl_175 br_175 wl_19 vdd gnd cell_6t
Xbit_r20_c175 bl_175 br_175 wl_20 vdd gnd cell_6t
Xbit_r21_c175 bl_175 br_175 wl_21 vdd gnd cell_6t
Xbit_r22_c175 bl_175 br_175 wl_22 vdd gnd cell_6t
Xbit_r23_c175 bl_175 br_175 wl_23 vdd gnd cell_6t
Xbit_r24_c175 bl_175 br_175 wl_24 vdd gnd cell_6t
Xbit_r25_c175 bl_175 br_175 wl_25 vdd gnd cell_6t
Xbit_r26_c175 bl_175 br_175 wl_26 vdd gnd cell_6t
Xbit_r27_c175 bl_175 br_175 wl_27 vdd gnd cell_6t
Xbit_r28_c175 bl_175 br_175 wl_28 vdd gnd cell_6t
Xbit_r29_c175 bl_175 br_175 wl_29 vdd gnd cell_6t
Xbit_r30_c175 bl_175 br_175 wl_30 vdd gnd cell_6t
Xbit_r31_c175 bl_175 br_175 wl_31 vdd gnd cell_6t
Xbit_r32_c175 bl_175 br_175 wl_32 vdd gnd cell_6t
Xbit_r33_c175 bl_175 br_175 wl_33 vdd gnd cell_6t
Xbit_r34_c175 bl_175 br_175 wl_34 vdd gnd cell_6t
Xbit_r35_c175 bl_175 br_175 wl_35 vdd gnd cell_6t
Xbit_r36_c175 bl_175 br_175 wl_36 vdd gnd cell_6t
Xbit_r37_c175 bl_175 br_175 wl_37 vdd gnd cell_6t
Xbit_r38_c175 bl_175 br_175 wl_38 vdd gnd cell_6t
Xbit_r39_c175 bl_175 br_175 wl_39 vdd gnd cell_6t
Xbit_r40_c175 bl_175 br_175 wl_40 vdd gnd cell_6t
Xbit_r41_c175 bl_175 br_175 wl_41 vdd gnd cell_6t
Xbit_r42_c175 bl_175 br_175 wl_42 vdd gnd cell_6t
Xbit_r43_c175 bl_175 br_175 wl_43 vdd gnd cell_6t
Xbit_r44_c175 bl_175 br_175 wl_44 vdd gnd cell_6t
Xbit_r45_c175 bl_175 br_175 wl_45 vdd gnd cell_6t
Xbit_r46_c175 bl_175 br_175 wl_46 vdd gnd cell_6t
Xbit_r47_c175 bl_175 br_175 wl_47 vdd gnd cell_6t
Xbit_r48_c175 bl_175 br_175 wl_48 vdd gnd cell_6t
Xbit_r49_c175 bl_175 br_175 wl_49 vdd gnd cell_6t
Xbit_r50_c175 bl_175 br_175 wl_50 vdd gnd cell_6t
Xbit_r51_c175 bl_175 br_175 wl_51 vdd gnd cell_6t
Xbit_r52_c175 bl_175 br_175 wl_52 vdd gnd cell_6t
Xbit_r53_c175 bl_175 br_175 wl_53 vdd gnd cell_6t
Xbit_r54_c175 bl_175 br_175 wl_54 vdd gnd cell_6t
Xbit_r55_c175 bl_175 br_175 wl_55 vdd gnd cell_6t
Xbit_r56_c175 bl_175 br_175 wl_56 vdd gnd cell_6t
Xbit_r57_c175 bl_175 br_175 wl_57 vdd gnd cell_6t
Xbit_r58_c175 bl_175 br_175 wl_58 vdd gnd cell_6t
Xbit_r59_c175 bl_175 br_175 wl_59 vdd gnd cell_6t
Xbit_r60_c175 bl_175 br_175 wl_60 vdd gnd cell_6t
Xbit_r61_c175 bl_175 br_175 wl_61 vdd gnd cell_6t
Xbit_r62_c175 bl_175 br_175 wl_62 vdd gnd cell_6t
Xbit_r63_c175 bl_175 br_175 wl_63 vdd gnd cell_6t
Xbit_r64_c175 bl_175 br_175 wl_64 vdd gnd cell_6t
Xbit_r65_c175 bl_175 br_175 wl_65 vdd gnd cell_6t
Xbit_r66_c175 bl_175 br_175 wl_66 vdd gnd cell_6t
Xbit_r67_c175 bl_175 br_175 wl_67 vdd gnd cell_6t
Xbit_r68_c175 bl_175 br_175 wl_68 vdd gnd cell_6t
Xbit_r69_c175 bl_175 br_175 wl_69 vdd gnd cell_6t
Xbit_r70_c175 bl_175 br_175 wl_70 vdd gnd cell_6t
Xbit_r71_c175 bl_175 br_175 wl_71 vdd gnd cell_6t
Xbit_r72_c175 bl_175 br_175 wl_72 vdd gnd cell_6t
Xbit_r73_c175 bl_175 br_175 wl_73 vdd gnd cell_6t
Xbit_r74_c175 bl_175 br_175 wl_74 vdd gnd cell_6t
Xbit_r75_c175 bl_175 br_175 wl_75 vdd gnd cell_6t
Xbit_r76_c175 bl_175 br_175 wl_76 vdd gnd cell_6t
Xbit_r77_c175 bl_175 br_175 wl_77 vdd gnd cell_6t
Xbit_r78_c175 bl_175 br_175 wl_78 vdd gnd cell_6t
Xbit_r79_c175 bl_175 br_175 wl_79 vdd gnd cell_6t
Xbit_r80_c175 bl_175 br_175 wl_80 vdd gnd cell_6t
Xbit_r81_c175 bl_175 br_175 wl_81 vdd gnd cell_6t
Xbit_r82_c175 bl_175 br_175 wl_82 vdd gnd cell_6t
Xbit_r83_c175 bl_175 br_175 wl_83 vdd gnd cell_6t
Xbit_r84_c175 bl_175 br_175 wl_84 vdd gnd cell_6t
Xbit_r85_c175 bl_175 br_175 wl_85 vdd gnd cell_6t
Xbit_r86_c175 bl_175 br_175 wl_86 vdd gnd cell_6t
Xbit_r87_c175 bl_175 br_175 wl_87 vdd gnd cell_6t
Xbit_r88_c175 bl_175 br_175 wl_88 vdd gnd cell_6t
Xbit_r89_c175 bl_175 br_175 wl_89 vdd gnd cell_6t
Xbit_r90_c175 bl_175 br_175 wl_90 vdd gnd cell_6t
Xbit_r91_c175 bl_175 br_175 wl_91 vdd gnd cell_6t
Xbit_r92_c175 bl_175 br_175 wl_92 vdd gnd cell_6t
Xbit_r93_c175 bl_175 br_175 wl_93 vdd gnd cell_6t
Xbit_r94_c175 bl_175 br_175 wl_94 vdd gnd cell_6t
Xbit_r95_c175 bl_175 br_175 wl_95 vdd gnd cell_6t
Xbit_r96_c175 bl_175 br_175 wl_96 vdd gnd cell_6t
Xbit_r97_c175 bl_175 br_175 wl_97 vdd gnd cell_6t
Xbit_r98_c175 bl_175 br_175 wl_98 vdd gnd cell_6t
Xbit_r99_c175 bl_175 br_175 wl_99 vdd gnd cell_6t
Xbit_r100_c175 bl_175 br_175 wl_100 vdd gnd cell_6t
Xbit_r101_c175 bl_175 br_175 wl_101 vdd gnd cell_6t
Xbit_r102_c175 bl_175 br_175 wl_102 vdd gnd cell_6t
Xbit_r103_c175 bl_175 br_175 wl_103 vdd gnd cell_6t
Xbit_r104_c175 bl_175 br_175 wl_104 vdd gnd cell_6t
Xbit_r105_c175 bl_175 br_175 wl_105 vdd gnd cell_6t
Xbit_r106_c175 bl_175 br_175 wl_106 vdd gnd cell_6t
Xbit_r107_c175 bl_175 br_175 wl_107 vdd gnd cell_6t
Xbit_r108_c175 bl_175 br_175 wl_108 vdd gnd cell_6t
Xbit_r109_c175 bl_175 br_175 wl_109 vdd gnd cell_6t
Xbit_r110_c175 bl_175 br_175 wl_110 vdd gnd cell_6t
Xbit_r111_c175 bl_175 br_175 wl_111 vdd gnd cell_6t
Xbit_r112_c175 bl_175 br_175 wl_112 vdd gnd cell_6t
Xbit_r113_c175 bl_175 br_175 wl_113 vdd gnd cell_6t
Xbit_r114_c175 bl_175 br_175 wl_114 vdd gnd cell_6t
Xbit_r115_c175 bl_175 br_175 wl_115 vdd gnd cell_6t
Xbit_r116_c175 bl_175 br_175 wl_116 vdd gnd cell_6t
Xbit_r117_c175 bl_175 br_175 wl_117 vdd gnd cell_6t
Xbit_r118_c175 bl_175 br_175 wl_118 vdd gnd cell_6t
Xbit_r119_c175 bl_175 br_175 wl_119 vdd gnd cell_6t
Xbit_r120_c175 bl_175 br_175 wl_120 vdd gnd cell_6t
Xbit_r121_c175 bl_175 br_175 wl_121 vdd gnd cell_6t
Xbit_r122_c175 bl_175 br_175 wl_122 vdd gnd cell_6t
Xbit_r123_c175 bl_175 br_175 wl_123 vdd gnd cell_6t
Xbit_r124_c175 bl_175 br_175 wl_124 vdd gnd cell_6t
Xbit_r125_c175 bl_175 br_175 wl_125 vdd gnd cell_6t
Xbit_r126_c175 bl_175 br_175 wl_126 vdd gnd cell_6t
Xbit_r127_c175 bl_175 br_175 wl_127 vdd gnd cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd cell_6t
Xbit_r1_c176 bl_176 br_176 wl_1 vdd gnd cell_6t
Xbit_r2_c176 bl_176 br_176 wl_2 vdd gnd cell_6t
Xbit_r3_c176 bl_176 br_176 wl_3 vdd gnd cell_6t
Xbit_r4_c176 bl_176 br_176 wl_4 vdd gnd cell_6t
Xbit_r5_c176 bl_176 br_176 wl_5 vdd gnd cell_6t
Xbit_r6_c176 bl_176 br_176 wl_6 vdd gnd cell_6t
Xbit_r7_c176 bl_176 br_176 wl_7 vdd gnd cell_6t
Xbit_r8_c176 bl_176 br_176 wl_8 vdd gnd cell_6t
Xbit_r9_c176 bl_176 br_176 wl_9 vdd gnd cell_6t
Xbit_r10_c176 bl_176 br_176 wl_10 vdd gnd cell_6t
Xbit_r11_c176 bl_176 br_176 wl_11 vdd gnd cell_6t
Xbit_r12_c176 bl_176 br_176 wl_12 vdd gnd cell_6t
Xbit_r13_c176 bl_176 br_176 wl_13 vdd gnd cell_6t
Xbit_r14_c176 bl_176 br_176 wl_14 vdd gnd cell_6t
Xbit_r15_c176 bl_176 br_176 wl_15 vdd gnd cell_6t
Xbit_r16_c176 bl_176 br_176 wl_16 vdd gnd cell_6t
Xbit_r17_c176 bl_176 br_176 wl_17 vdd gnd cell_6t
Xbit_r18_c176 bl_176 br_176 wl_18 vdd gnd cell_6t
Xbit_r19_c176 bl_176 br_176 wl_19 vdd gnd cell_6t
Xbit_r20_c176 bl_176 br_176 wl_20 vdd gnd cell_6t
Xbit_r21_c176 bl_176 br_176 wl_21 vdd gnd cell_6t
Xbit_r22_c176 bl_176 br_176 wl_22 vdd gnd cell_6t
Xbit_r23_c176 bl_176 br_176 wl_23 vdd gnd cell_6t
Xbit_r24_c176 bl_176 br_176 wl_24 vdd gnd cell_6t
Xbit_r25_c176 bl_176 br_176 wl_25 vdd gnd cell_6t
Xbit_r26_c176 bl_176 br_176 wl_26 vdd gnd cell_6t
Xbit_r27_c176 bl_176 br_176 wl_27 vdd gnd cell_6t
Xbit_r28_c176 bl_176 br_176 wl_28 vdd gnd cell_6t
Xbit_r29_c176 bl_176 br_176 wl_29 vdd gnd cell_6t
Xbit_r30_c176 bl_176 br_176 wl_30 vdd gnd cell_6t
Xbit_r31_c176 bl_176 br_176 wl_31 vdd gnd cell_6t
Xbit_r32_c176 bl_176 br_176 wl_32 vdd gnd cell_6t
Xbit_r33_c176 bl_176 br_176 wl_33 vdd gnd cell_6t
Xbit_r34_c176 bl_176 br_176 wl_34 vdd gnd cell_6t
Xbit_r35_c176 bl_176 br_176 wl_35 vdd gnd cell_6t
Xbit_r36_c176 bl_176 br_176 wl_36 vdd gnd cell_6t
Xbit_r37_c176 bl_176 br_176 wl_37 vdd gnd cell_6t
Xbit_r38_c176 bl_176 br_176 wl_38 vdd gnd cell_6t
Xbit_r39_c176 bl_176 br_176 wl_39 vdd gnd cell_6t
Xbit_r40_c176 bl_176 br_176 wl_40 vdd gnd cell_6t
Xbit_r41_c176 bl_176 br_176 wl_41 vdd gnd cell_6t
Xbit_r42_c176 bl_176 br_176 wl_42 vdd gnd cell_6t
Xbit_r43_c176 bl_176 br_176 wl_43 vdd gnd cell_6t
Xbit_r44_c176 bl_176 br_176 wl_44 vdd gnd cell_6t
Xbit_r45_c176 bl_176 br_176 wl_45 vdd gnd cell_6t
Xbit_r46_c176 bl_176 br_176 wl_46 vdd gnd cell_6t
Xbit_r47_c176 bl_176 br_176 wl_47 vdd gnd cell_6t
Xbit_r48_c176 bl_176 br_176 wl_48 vdd gnd cell_6t
Xbit_r49_c176 bl_176 br_176 wl_49 vdd gnd cell_6t
Xbit_r50_c176 bl_176 br_176 wl_50 vdd gnd cell_6t
Xbit_r51_c176 bl_176 br_176 wl_51 vdd gnd cell_6t
Xbit_r52_c176 bl_176 br_176 wl_52 vdd gnd cell_6t
Xbit_r53_c176 bl_176 br_176 wl_53 vdd gnd cell_6t
Xbit_r54_c176 bl_176 br_176 wl_54 vdd gnd cell_6t
Xbit_r55_c176 bl_176 br_176 wl_55 vdd gnd cell_6t
Xbit_r56_c176 bl_176 br_176 wl_56 vdd gnd cell_6t
Xbit_r57_c176 bl_176 br_176 wl_57 vdd gnd cell_6t
Xbit_r58_c176 bl_176 br_176 wl_58 vdd gnd cell_6t
Xbit_r59_c176 bl_176 br_176 wl_59 vdd gnd cell_6t
Xbit_r60_c176 bl_176 br_176 wl_60 vdd gnd cell_6t
Xbit_r61_c176 bl_176 br_176 wl_61 vdd gnd cell_6t
Xbit_r62_c176 bl_176 br_176 wl_62 vdd gnd cell_6t
Xbit_r63_c176 bl_176 br_176 wl_63 vdd gnd cell_6t
Xbit_r64_c176 bl_176 br_176 wl_64 vdd gnd cell_6t
Xbit_r65_c176 bl_176 br_176 wl_65 vdd gnd cell_6t
Xbit_r66_c176 bl_176 br_176 wl_66 vdd gnd cell_6t
Xbit_r67_c176 bl_176 br_176 wl_67 vdd gnd cell_6t
Xbit_r68_c176 bl_176 br_176 wl_68 vdd gnd cell_6t
Xbit_r69_c176 bl_176 br_176 wl_69 vdd gnd cell_6t
Xbit_r70_c176 bl_176 br_176 wl_70 vdd gnd cell_6t
Xbit_r71_c176 bl_176 br_176 wl_71 vdd gnd cell_6t
Xbit_r72_c176 bl_176 br_176 wl_72 vdd gnd cell_6t
Xbit_r73_c176 bl_176 br_176 wl_73 vdd gnd cell_6t
Xbit_r74_c176 bl_176 br_176 wl_74 vdd gnd cell_6t
Xbit_r75_c176 bl_176 br_176 wl_75 vdd gnd cell_6t
Xbit_r76_c176 bl_176 br_176 wl_76 vdd gnd cell_6t
Xbit_r77_c176 bl_176 br_176 wl_77 vdd gnd cell_6t
Xbit_r78_c176 bl_176 br_176 wl_78 vdd gnd cell_6t
Xbit_r79_c176 bl_176 br_176 wl_79 vdd gnd cell_6t
Xbit_r80_c176 bl_176 br_176 wl_80 vdd gnd cell_6t
Xbit_r81_c176 bl_176 br_176 wl_81 vdd gnd cell_6t
Xbit_r82_c176 bl_176 br_176 wl_82 vdd gnd cell_6t
Xbit_r83_c176 bl_176 br_176 wl_83 vdd gnd cell_6t
Xbit_r84_c176 bl_176 br_176 wl_84 vdd gnd cell_6t
Xbit_r85_c176 bl_176 br_176 wl_85 vdd gnd cell_6t
Xbit_r86_c176 bl_176 br_176 wl_86 vdd gnd cell_6t
Xbit_r87_c176 bl_176 br_176 wl_87 vdd gnd cell_6t
Xbit_r88_c176 bl_176 br_176 wl_88 vdd gnd cell_6t
Xbit_r89_c176 bl_176 br_176 wl_89 vdd gnd cell_6t
Xbit_r90_c176 bl_176 br_176 wl_90 vdd gnd cell_6t
Xbit_r91_c176 bl_176 br_176 wl_91 vdd gnd cell_6t
Xbit_r92_c176 bl_176 br_176 wl_92 vdd gnd cell_6t
Xbit_r93_c176 bl_176 br_176 wl_93 vdd gnd cell_6t
Xbit_r94_c176 bl_176 br_176 wl_94 vdd gnd cell_6t
Xbit_r95_c176 bl_176 br_176 wl_95 vdd gnd cell_6t
Xbit_r96_c176 bl_176 br_176 wl_96 vdd gnd cell_6t
Xbit_r97_c176 bl_176 br_176 wl_97 vdd gnd cell_6t
Xbit_r98_c176 bl_176 br_176 wl_98 vdd gnd cell_6t
Xbit_r99_c176 bl_176 br_176 wl_99 vdd gnd cell_6t
Xbit_r100_c176 bl_176 br_176 wl_100 vdd gnd cell_6t
Xbit_r101_c176 bl_176 br_176 wl_101 vdd gnd cell_6t
Xbit_r102_c176 bl_176 br_176 wl_102 vdd gnd cell_6t
Xbit_r103_c176 bl_176 br_176 wl_103 vdd gnd cell_6t
Xbit_r104_c176 bl_176 br_176 wl_104 vdd gnd cell_6t
Xbit_r105_c176 bl_176 br_176 wl_105 vdd gnd cell_6t
Xbit_r106_c176 bl_176 br_176 wl_106 vdd gnd cell_6t
Xbit_r107_c176 bl_176 br_176 wl_107 vdd gnd cell_6t
Xbit_r108_c176 bl_176 br_176 wl_108 vdd gnd cell_6t
Xbit_r109_c176 bl_176 br_176 wl_109 vdd gnd cell_6t
Xbit_r110_c176 bl_176 br_176 wl_110 vdd gnd cell_6t
Xbit_r111_c176 bl_176 br_176 wl_111 vdd gnd cell_6t
Xbit_r112_c176 bl_176 br_176 wl_112 vdd gnd cell_6t
Xbit_r113_c176 bl_176 br_176 wl_113 vdd gnd cell_6t
Xbit_r114_c176 bl_176 br_176 wl_114 vdd gnd cell_6t
Xbit_r115_c176 bl_176 br_176 wl_115 vdd gnd cell_6t
Xbit_r116_c176 bl_176 br_176 wl_116 vdd gnd cell_6t
Xbit_r117_c176 bl_176 br_176 wl_117 vdd gnd cell_6t
Xbit_r118_c176 bl_176 br_176 wl_118 vdd gnd cell_6t
Xbit_r119_c176 bl_176 br_176 wl_119 vdd gnd cell_6t
Xbit_r120_c176 bl_176 br_176 wl_120 vdd gnd cell_6t
Xbit_r121_c176 bl_176 br_176 wl_121 vdd gnd cell_6t
Xbit_r122_c176 bl_176 br_176 wl_122 vdd gnd cell_6t
Xbit_r123_c176 bl_176 br_176 wl_123 vdd gnd cell_6t
Xbit_r124_c176 bl_176 br_176 wl_124 vdd gnd cell_6t
Xbit_r125_c176 bl_176 br_176 wl_125 vdd gnd cell_6t
Xbit_r126_c176 bl_176 br_176 wl_126 vdd gnd cell_6t
Xbit_r127_c176 bl_176 br_176 wl_127 vdd gnd cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd cell_6t
Xbit_r1_c177 bl_177 br_177 wl_1 vdd gnd cell_6t
Xbit_r2_c177 bl_177 br_177 wl_2 vdd gnd cell_6t
Xbit_r3_c177 bl_177 br_177 wl_3 vdd gnd cell_6t
Xbit_r4_c177 bl_177 br_177 wl_4 vdd gnd cell_6t
Xbit_r5_c177 bl_177 br_177 wl_5 vdd gnd cell_6t
Xbit_r6_c177 bl_177 br_177 wl_6 vdd gnd cell_6t
Xbit_r7_c177 bl_177 br_177 wl_7 vdd gnd cell_6t
Xbit_r8_c177 bl_177 br_177 wl_8 vdd gnd cell_6t
Xbit_r9_c177 bl_177 br_177 wl_9 vdd gnd cell_6t
Xbit_r10_c177 bl_177 br_177 wl_10 vdd gnd cell_6t
Xbit_r11_c177 bl_177 br_177 wl_11 vdd gnd cell_6t
Xbit_r12_c177 bl_177 br_177 wl_12 vdd gnd cell_6t
Xbit_r13_c177 bl_177 br_177 wl_13 vdd gnd cell_6t
Xbit_r14_c177 bl_177 br_177 wl_14 vdd gnd cell_6t
Xbit_r15_c177 bl_177 br_177 wl_15 vdd gnd cell_6t
Xbit_r16_c177 bl_177 br_177 wl_16 vdd gnd cell_6t
Xbit_r17_c177 bl_177 br_177 wl_17 vdd gnd cell_6t
Xbit_r18_c177 bl_177 br_177 wl_18 vdd gnd cell_6t
Xbit_r19_c177 bl_177 br_177 wl_19 vdd gnd cell_6t
Xbit_r20_c177 bl_177 br_177 wl_20 vdd gnd cell_6t
Xbit_r21_c177 bl_177 br_177 wl_21 vdd gnd cell_6t
Xbit_r22_c177 bl_177 br_177 wl_22 vdd gnd cell_6t
Xbit_r23_c177 bl_177 br_177 wl_23 vdd gnd cell_6t
Xbit_r24_c177 bl_177 br_177 wl_24 vdd gnd cell_6t
Xbit_r25_c177 bl_177 br_177 wl_25 vdd gnd cell_6t
Xbit_r26_c177 bl_177 br_177 wl_26 vdd gnd cell_6t
Xbit_r27_c177 bl_177 br_177 wl_27 vdd gnd cell_6t
Xbit_r28_c177 bl_177 br_177 wl_28 vdd gnd cell_6t
Xbit_r29_c177 bl_177 br_177 wl_29 vdd gnd cell_6t
Xbit_r30_c177 bl_177 br_177 wl_30 vdd gnd cell_6t
Xbit_r31_c177 bl_177 br_177 wl_31 vdd gnd cell_6t
Xbit_r32_c177 bl_177 br_177 wl_32 vdd gnd cell_6t
Xbit_r33_c177 bl_177 br_177 wl_33 vdd gnd cell_6t
Xbit_r34_c177 bl_177 br_177 wl_34 vdd gnd cell_6t
Xbit_r35_c177 bl_177 br_177 wl_35 vdd gnd cell_6t
Xbit_r36_c177 bl_177 br_177 wl_36 vdd gnd cell_6t
Xbit_r37_c177 bl_177 br_177 wl_37 vdd gnd cell_6t
Xbit_r38_c177 bl_177 br_177 wl_38 vdd gnd cell_6t
Xbit_r39_c177 bl_177 br_177 wl_39 vdd gnd cell_6t
Xbit_r40_c177 bl_177 br_177 wl_40 vdd gnd cell_6t
Xbit_r41_c177 bl_177 br_177 wl_41 vdd gnd cell_6t
Xbit_r42_c177 bl_177 br_177 wl_42 vdd gnd cell_6t
Xbit_r43_c177 bl_177 br_177 wl_43 vdd gnd cell_6t
Xbit_r44_c177 bl_177 br_177 wl_44 vdd gnd cell_6t
Xbit_r45_c177 bl_177 br_177 wl_45 vdd gnd cell_6t
Xbit_r46_c177 bl_177 br_177 wl_46 vdd gnd cell_6t
Xbit_r47_c177 bl_177 br_177 wl_47 vdd gnd cell_6t
Xbit_r48_c177 bl_177 br_177 wl_48 vdd gnd cell_6t
Xbit_r49_c177 bl_177 br_177 wl_49 vdd gnd cell_6t
Xbit_r50_c177 bl_177 br_177 wl_50 vdd gnd cell_6t
Xbit_r51_c177 bl_177 br_177 wl_51 vdd gnd cell_6t
Xbit_r52_c177 bl_177 br_177 wl_52 vdd gnd cell_6t
Xbit_r53_c177 bl_177 br_177 wl_53 vdd gnd cell_6t
Xbit_r54_c177 bl_177 br_177 wl_54 vdd gnd cell_6t
Xbit_r55_c177 bl_177 br_177 wl_55 vdd gnd cell_6t
Xbit_r56_c177 bl_177 br_177 wl_56 vdd gnd cell_6t
Xbit_r57_c177 bl_177 br_177 wl_57 vdd gnd cell_6t
Xbit_r58_c177 bl_177 br_177 wl_58 vdd gnd cell_6t
Xbit_r59_c177 bl_177 br_177 wl_59 vdd gnd cell_6t
Xbit_r60_c177 bl_177 br_177 wl_60 vdd gnd cell_6t
Xbit_r61_c177 bl_177 br_177 wl_61 vdd gnd cell_6t
Xbit_r62_c177 bl_177 br_177 wl_62 vdd gnd cell_6t
Xbit_r63_c177 bl_177 br_177 wl_63 vdd gnd cell_6t
Xbit_r64_c177 bl_177 br_177 wl_64 vdd gnd cell_6t
Xbit_r65_c177 bl_177 br_177 wl_65 vdd gnd cell_6t
Xbit_r66_c177 bl_177 br_177 wl_66 vdd gnd cell_6t
Xbit_r67_c177 bl_177 br_177 wl_67 vdd gnd cell_6t
Xbit_r68_c177 bl_177 br_177 wl_68 vdd gnd cell_6t
Xbit_r69_c177 bl_177 br_177 wl_69 vdd gnd cell_6t
Xbit_r70_c177 bl_177 br_177 wl_70 vdd gnd cell_6t
Xbit_r71_c177 bl_177 br_177 wl_71 vdd gnd cell_6t
Xbit_r72_c177 bl_177 br_177 wl_72 vdd gnd cell_6t
Xbit_r73_c177 bl_177 br_177 wl_73 vdd gnd cell_6t
Xbit_r74_c177 bl_177 br_177 wl_74 vdd gnd cell_6t
Xbit_r75_c177 bl_177 br_177 wl_75 vdd gnd cell_6t
Xbit_r76_c177 bl_177 br_177 wl_76 vdd gnd cell_6t
Xbit_r77_c177 bl_177 br_177 wl_77 vdd gnd cell_6t
Xbit_r78_c177 bl_177 br_177 wl_78 vdd gnd cell_6t
Xbit_r79_c177 bl_177 br_177 wl_79 vdd gnd cell_6t
Xbit_r80_c177 bl_177 br_177 wl_80 vdd gnd cell_6t
Xbit_r81_c177 bl_177 br_177 wl_81 vdd gnd cell_6t
Xbit_r82_c177 bl_177 br_177 wl_82 vdd gnd cell_6t
Xbit_r83_c177 bl_177 br_177 wl_83 vdd gnd cell_6t
Xbit_r84_c177 bl_177 br_177 wl_84 vdd gnd cell_6t
Xbit_r85_c177 bl_177 br_177 wl_85 vdd gnd cell_6t
Xbit_r86_c177 bl_177 br_177 wl_86 vdd gnd cell_6t
Xbit_r87_c177 bl_177 br_177 wl_87 vdd gnd cell_6t
Xbit_r88_c177 bl_177 br_177 wl_88 vdd gnd cell_6t
Xbit_r89_c177 bl_177 br_177 wl_89 vdd gnd cell_6t
Xbit_r90_c177 bl_177 br_177 wl_90 vdd gnd cell_6t
Xbit_r91_c177 bl_177 br_177 wl_91 vdd gnd cell_6t
Xbit_r92_c177 bl_177 br_177 wl_92 vdd gnd cell_6t
Xbit_r93_c177 bl_177 br_177 wl_93 vdd gnd cell_6t
Xbit_r94_c177 bl_177 br_177 wl_94 vdd gnd cell_6t
Xbit_r95_c177 bl_177 br_177 wl_95 vdd gnd cell_6t
Xbit_r96_c177 bl_177 br_177 wl_96 vdd gnd cell_6t
Xbit_r97_c177 bl_177 br_177 wl_97 vdd gnd cell_6t
Xbit_r98_c177 bl_177 br_177 wl_98 vdd gnd cell_6t
Xbit_r99_c177 bl_177 br_177 wl_99 vdd gnd cell_6t
Xbit_r100_c177 bl_177 br_177 wl_100 vdd gnd cell_6t
Xbit_r101_c177 bl_177 br_177 wl_101 vdd gnd cell_6t
Xbit_r102_c177 bl_177 br_177 wl_102 vdd gnd cell_6t
Xbit_r103_c177 bl_177 br_177 wl_103 vdd gnd cell_6t
Xbit_r104_c177 bl_177 br_177 wl_104 vdd gnd cell_6t
Xbit_r105_c177 bl_177 br_177 wl_105 vdd gnd cell_6t
Xbit_r106_c177 bl_177 br_177 wl_106 vdd gnd cell_6t
Xbit_r107_c177 bl_177 br_177 wl_107 vdd gnd cell_6t
Xbit_r108_c177 bl_177 br_177 wl_108 vdd gnd cell_6t
Xbit_r109_c177 bl_177 br_177 wl_109 vdd gnd cell_6t
Xbit_r110_c177 bl_177 br_177 wl_110 vdd gnd cell_6t
Xbit_r111_c177 bl_177 br_177 wl_111 vdd gnd cell_6t
Xbit_r112_c177 bl_177 br_177 wl_112 vdd gnd cell_6t
Xbit_r113_c177 bl_177 br_177 wl_113 vdd gnd cell_6t
Xbit_r114_c177 bl_177 br_177 wl_114 vdd gnd cell_6t
Xbit_r115_c177 bl_177 br_177 wl_115 vdd gnd cell_6t
Xbit_r116_c177 bl_177 br_177 wl_116 vdd gnd cell_6t
Xbit_r117_c177 bl_177 br_177 wl_117 vdd gnd cell_6t
Xbit_r118_c177 bl_177 br_177 wl_118 vdd gnd cell_6t
Xbit_r119_c177 bl_177 br_177 wl_119 vdd gnd cell_6t
Xbit_r120_c177 bl_177 br_177 wl_120 vdd gnd cell_6t
Xbit_r121_c177 bl_177 br_177 wl_121 vdd gnd cell_6t
Xbit_r122_c177 bl_177 br_177 wl_122 vdd gnd cell_6t
Xbit_r123_c177 bl_177 br_177 wl_123 vdd gnd cell_6t
Xbit_r124_c177 bl_177 br_177 wl_124 vdd gnd cell_6t
Xbit_r125_c177 bl_177 br_177 wl_125 vdd gnd cell_6t
Xbit_r126_c177 bl_177 br_177 wl_126 vdd gnd cell_6t
Xbit_r127_c177 bl_177 br_177 wl_127 vdd gnd cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd cell_6t
Xbit_r1_c178 bl_178 br_178 wl_1 vdd gnd cell_6t
Xbit_r2_c178 bl_178 br_178 wl_2 vdd gnd cell_6t
Xbit_r3_c178 bl_178 br_178 wl_3 vdd gnd cell_6t
Xbit_r4_c178 bl_178 br_178 wl_4 vdd gnd cell_6t
Xbit_r5_c178 bl_178 br_178 wl_5 vdd gnd cell_6t
Xbit_r6_c178 bl_178 br_178 wl_6 vdd gnd cell_6t
Xbit_r7_c178 bl_178 br_178 wl_7 vdd gnd cell_6t
Xbit_r8_c178 bl_178 br_178 wl_8 vdd gnd cell_6t
Xbit_r9_c178 bl_178 br_178 wl_9 vdd gnd cell_6t
Xbit_r10_c178 bl_178 br_178 wl_10 vdd gnd cell_6t
Xbit_r11_c178 bl_178 br_178 wl_11 vdd gnd cell_6t
Xbit_r12_c178 bl_178 br_178 wl_12 vdd gnd cell_6t
Xbit_r13_c178 bl_178 br_178 wl_13 vdd gnd cell_6t
Xbit_r14_c178 bl_178 br_178 wl_14 vdd gnd cell_6t
Xbit_r15_c178 bl_178 br_178 wl_15 vdd gnd cell_6t
Xbit_r16_c178 bl_178 br_178 wl_16 vdd gnd cell_6t
Xbit_r17_c178 bl_178 br_178 wl_17 vdd gnd cell_6t
Xbit_r18_c178 bl_178 br_178 wl_18 vdd gnd cell_6t
Xbit_r19_c178 bl_178 br_178 wl_19 vdd gnd cell_6t
Xbit_r20_c178 bl_178 br_178 wl_20 vdd gnd cell_6t
Xbit_r21_c178 bl_178 br_178 wl_21 vdd gnd cell_6t
Xbit_r22_c178 bl_178 br_178 wl_22 vdd gnd cell_6t
Xbit_r23_c178 bl_178 br_178 wl_23 vdd gnd cell_6t
Xbit_r24_c178 bl_178 br_178 wl_24 vdd gnd cell_6t
Xbit_r25_c178 bl_178 br_178 wl_25 vdd gnd cell_6t
Xbit_r26_c178 bl_178 br_178 wl_26 vdd gnd cell_6t
Xbit_r27_c178 bl_178 br_178 wl_27 vdd gnd cell_6t
Xbit_r28_c178 bl_178 br_178 wl_28 vdd gnd cell_6t
Xbit_r29_c178 bl_178 br_178 wl_29 vdd gnd cell_6t
Xbit_r30_c178 bl_178 br_178 wl_30 vdd gnd cell_6t
Xbit_r31_c178 bl_178 br_178 wl_31 vdd gnd cell_6t
Xbit_r32_c178 bl_178 br_178 wl_32 vdd gnd cell_6t
Xbit_r33_c178 bl_178 br_178 wl_33 vdd gnd cell_6t
Xbit_r34_c178 bl_178 br_178 wl_34 vdd gnd cell_6t
Xbit_r35_c178 bl_178 br_178 wl_35 vdd gnd cell_6t
Xbit_r36_c178 bl_178 br_178 wl_36 vdd gnd cell_6t
Xbit_r37_c178 bl_178 br_178 wl_37 vdd gnd cell_6t
Xbit_r38_c178 bl_178 br_178 wl_38 vdd gnd cell_6t
Xbit_r39_c178 bl_178 br_178 wl_39 vdd gnd cell_6t
Xbit_r40_c178 bl_178 br_178 wl_40 vdd gnd cell_6t
Xbit_r41_c178 bl_178 br_178 wl_41 vdd gnd cell_6t
Xbit_r42_c178 bl_178 br_178 wl_42 vdd gnd cell_6t
Xbit_r43_c178 bl_178 br_178 wl_43 vdd gnd cell_6t
Xbit_r44_c178 bl_178 br_178 wl_44 vdd gnd cell_6t
Xbit_r45_c178 bl_178 br_178 wl_45 vdd gnd cell_6t
Xbit_r46_c178 bl_178 br_178 wl_46 vdd gnd cell_6t
Xbit_r47_c178 bl_178 br_178 wl_47 vdd gnd cell_6t
Xbit_r48_c178 bl_178 br_178 wl_48 vdd gnd cell_6t
Xbit_r49_c178 bl_178 br_178 wl_49 vdd gnd cell_6t
Xbit_r50_c178 bl_178 br_178 wl_50 vdd gnd cell_6t
Xbit_r51_c178 bl_178 br_178 wl_51 vdd gnd cell_6t
Xbit_r52_c178 bl_178 br_178 wl_52 vdd gnd cell_6t
Xbit_r53_c178 bl_178 br_178 wl_53 vdd gnd cell_6t
Xbit_r54_c178 bl_178 br_178 wl_54 vdd gnd cell_6t
Xbit_r55_c178 bl_178 br_178 wl_55 vdd gnd cell_6t
Xbit_r56_c178 bl_178 br_178 wl_56 vdd gnd cell_6t
Xbit_r57_c178 bl_178 br_178 wl_57 vdd gnd cell_6t
Xbit_r58_c178 bl_178 br_178 wl_58 vdd gnd cell_6t
Xbit_r59_c178 bl_178 br_178 wl_59 vdd gnd cell_6t
Xbit_r60_c178 bl_178 br_178 wl_60 vdd gnd cell_6t
Xbit_r61_c178 bl_178 br_178 wl_61 vdd gnd cell_6t
Xbit_r62_c178 bl_178 br_178 wl_62 vdd gnd cell_6t
Xbit_r63_c178 bl_178 br_178 wl_63 vdd gnd cell_6t
Xbit_r64_c178 bl_178 br_178 wl_64 vdd gnd cell_6t
Xbit_r65_c178 bl_178 br_178 wl_65 vdd gnd cell_6t
Xbit_r66_c178 bl_178 br_178 wl_66 vdd gnd cell_6t
Xbit_r67_c178 bl_178 br_178 wl_67 vdd gnd cell_6t
Xbit_r68_c178 bl_178 br_178 wl_68 vdd gnd cell_6t
Xbit_r69_c178 bl_178 br_178 wl_69 vdd gnd cell_6t
Xbit_r70_c178 bl_178 br_178 wl_70 vdd gnd cell_6t
Xbit_r71_c178 bl_178 br_178 wl_71 vdd gnd cell_6t
Xbit_r72_c178 bl_178 br_178 wl_72 vdd gnd cell_6t
Xbit_r73_c178 bl_178 br_178 wl_73 vdd gnd cell_6t
Xbit_r74_c178 bl_178 br_178 wl_74 vdd gnd cell_6t
Xbit_r75_c178 bl_178 br_178 wl_75 vdd gnd cell_6t
Xbit_r76_c178 bl_178 br_178 wl_76 vdd gnd cell_6t
Xbit_r77_c178 bl_178 br_178 wl_77 vdd gnd cell_6t
Xbit_r78_c178 bl_178 br_178 wl_78 vdd gnd cell_6t
Xbit_r79_c178 bl_178 br_178 wl_79 vdd gnd cell_6t
Xbit_r80_c178 bl_178 br_178 wl_80 vdd gnd cell_6t
Xbit_r81_c178 bl_178 br_178 wl_81 vdd gnd cell_6t
Xbit_r82_c178 bl_178 br_178 wl_82 vdd gnd cell_6t
Xbit_r83_c178 bl_178 br_178 wl_83 vdd gnd cell_6t
Xbit_r84_c178 bl_178 br_178 wl_84 vdd gnd cell_6t
Xbit_r85_c178 bl_178 br_178 wl_85 vdd gnd cell_6t
Xbit_r86_c178 bl_178 br_178 wl_86 vdd gnd cell_6t
Xbit_r87_c178 bl_178 br_178 wl_87 vdd gnd cell_6t
Xbit_r88_c178 bl_178 br_178 wl_88 vdd gnd cell_6t
Xbit_r89_c178 bl_178 br_178 wl_89 vdd gnd cell_6t
Xbit_r90_c178 bl_178 br_178 wl_90 vdd gnd cell_6t
Xbit_r91_c178 bl_178 br_178 wl_91 vdd gnd cell_6t
Xbit_r92_c178 bl_178 br_178 wl_92 vdd gnd cell_6t
Xbit_r93_c178 bl_178 br_178 wl_93 vdd gnd cell_6t
Xbit_r94_c178 bl_178 br_178 wl_94 vdd gnd cell_6t
Xbit_r95_c178 bl_178 br_178 wl_95 vdd gnd cell_6t
Xbit_r96_c178 bl_178 br_178 wl_96 vdd gnd cell_6t
Xbit_r97_c178 bl_178 br_178 wl_97 vdd gnd cell_6t
Xbit_r98_c178 bl_178 br_178 wl_98 vdd gnd cell_6t
Xbit_r99_c178 bl_178 br_178 wl_99 vdd gnd cell_6t
Xbit_r100_c178 bl_178 br_178 wl_100 vdd gnd cell_6t
Xbit_r101_c178 bl_178 br_178 wl_101 vdd gnd cell_6t
Xbit_r102_c178 bl_178 br_178 wl_102 vdd gnd cell_6t
Xbit_r103_c178 bl_178 br_178 wl_103 vdd gnd cell_6t
Xbit_r104_c178 bl_178 br_178 wl_104 vdd gnd cell_6t
Xbit_r105_c178 bl_178 br_178 wl_105 vdd gnd cell_6t
Xbit_r106_c178 bl_178 br_178 wl_106 vdd gnd cell_6t
Xbit_r107_c178 bl_178 br_178 wl_107 vdd gnd cell_6t
Xbit_r108_c178 bl_178 br_178 wl_108 vdd gnd cell_6t
Xbit_r109_c178 bl_178 br_178 wl_109 vdd gnd cell_6t
Xbit_r110_c178 bl_178 br_178 wl_110 vdd gnd cell_6t
Xbit_r111_c178 bl_178 br_178 wl_111 vdd gnd cell_6t
Xbit_r112_c178 bl_178 br_178 wl_112 vdd gnd cell_6t
Xbit_r113_c178 bl_178 br_178 wl_113 vdd gnd cell_6t
Xbit_r114_c178 bl_178 br_178 wl_114 vdd gnd cell_6t
Xbit_r115_c178 bl_178 br_178 wl_115 vdd gnd cell_6t
Xbit_r116_c178 bl_178 br_178 wl_116 vdd gnd cell_6t
Xbit_r117_c178 bl_178 br_178 wl_117 vdd gnd cell_6t
Xbit_r118_c178 bl_178 br_178 wl_118 vdd gnd cell_6t
Xbit_r119_c178 bl_178 br_178 wl_119 vdd gnd cell_6t
Xbit_r120_c178 bl_178 br_178 wl_120 vdd gnd cell_6t
Xbit_r121_c178 bl_178 br_178 wl_121 vdd gnd cell_6t
Xbit_r122_c178 bl_178 br_178 wl_122 vdd gnd cell_6t
Xbit_r123_c178 bl_178 br_178 wl_123 vdd gnd cell_6t
Xbit_r124_c178 bl_178 br_178 wl_124 vdd gnd cell_6t
Xbit_r125_c178 bl_178 br_178 wl_125 vdd gnd cell_6t
Xbit_r126_c178 bl_178 br_178 wl_126 vdd gnd cell_6t
Xbit_r127_c178 bl_178 br_178 wl_127 vdd gnd cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd cell_6t
Xbit_r1_c179 bl_179 br_179 wl_1 vdd gnd cell_6t
Xbit_r2_c179 bl_179 br_179 wl_2 vdd gnd cell_6t
Xbit_r3_c179 bl_179 br_179 wl_3 vdd gnd cell_6t
Xbit_r4_c179 bl_179 br_179 wl_4 vdd gnd cell_6t
Xbit_r5_c179 bl_179 br_179 wl_5 vdd gnd cell_6t
Xbit_r6_c179 bl_179 br_179 wl_6 vdd gnd cell_6t
Xbit_r7_c179 bl_179 br_179 wl_7 vdd gnd cell_6t
Xbit_r8_c179 bl_179 br_179 wl_8 vdd gnd cell_6t
Xbit_r9_c179 bl_179 br_179 wl_9 vdd gnd cell_6t
Xbit_r10_c179 bl_179 br_179 wl_10 vdd gnd cell_6t
Xbit_r11_c179 bl_179 br_179 wl_11 vdd gnd cell_6t
Xbit_r12_c179 bl_179 br_179 wl_12 vdd gnd cell_6t
Xbit_r13_c179 bl_179 br_179 wl_13 vdd gnd cell_6t
Xbit_r14_c179 bl_179 br_179 wl_14 vdd gnd cell_6t
Xbit_r15_c179 bl_179 br_179 wl_15 vdd gnd cell_6t
Xbit_r16_c179 bl_179 br_179 wl_16 vdd gnd cell_6t
Xbit_r17_c179 bl_179 br_179 wl_17 vdd gnd cell_6t
Xbit_r18_c179 bl_179 br_179 wl_18 vdd gnd cell_6t
Xbit_r19_c179 bl_179 br_179 wl_19 vdd gnd cell_6t
Xbit_r20_c179 bl_179 br_179 wl_20 vdd gnd cell_6t
Xbit_r21_c179 bl_179 br_179 wl_21 vdd gnd cell_6t
Xbit_r22_c179 bl_179 br_179 wl_22 vdd gnd cell_6t
Xbit_r23_c179 bl_179 br_179 wl_23 vdd gnd cell_6t
Xbit_r24_c179 bl_179 br_179 wl_24 vdd gnd cell_6t
Xbit_r25_c179 bl_179 br_179 wl_25 vdd gnd cell_6t
Xbit_r26_c179 bl_179 br_179 wl_26 vdd gnd cell_6t
Xbit_r27_c179 bl_179 br_179 wl_27 vdd gnd cell_6t
Xbit_r28_c179 bl_179 br_179 wl_28 vdd gnd cell_6t
Xbit_r29_c179 bl_179 br_179 wl_29 vdd gnd cell_6t
Xbit_r30_c179 bl_179 br_179 wl_30 vdd gnd cell_6t
Xbit_r31_c179 bl_179 br_179 wl_31 vdd gnd cell_6t
Xbit_r32_c179 bl_179 br_179 wl_32 vdd gnd cell_6t
Xbit_r33_c179 bl_179 br_179 wl_33 vdd gnd cell_6t
Xbit_r34_c179 bl_179 br_179 wl_34 vdd gnd cell_6t
Xbit_r35_c179 bl_179 br_179 wl_35 vdd gnd cell_6t
Xbit_r36_c179 bl_179 br_179 wl_36 vdd gnd cell_6t
Xbit_r37_c179 bl_179 br_179 wl_37 vdd gnd cell_6t
Xbit_r38_c179 bl_179 br_179 wl_38 vdd gnd cell_6t
Xbit_r39_c179 bl_179 br_179 wl_39 vdd gnd cell_6t
Xbit_r40_c179 bl_179 br_179 wl_40 vdd gnd cell_6t
Xbit_r41_c179 bl_179 br_179 wl_41 vdd gnd cell_6t
Xbit_r42_c179 bl_179 br_179 wl_42 vdd gnd cell_6t
Xbit_r43_c179 bl_179 br_179 wl_43 vdd gnd cell_6t
Xbit_r44_c179 bl_179 br_179 wl_44 vdd gnd cell_6t
Xbit_r45_c179 bl_179 br_179 wl_45 vdd gnd cell_6t
Xbit_r46_c179 bl_179 br_179 wl_46 vdd gnd cell_6t
Xbit_r47_c179 bl_179 br_179 wl_47 vdd gnd cell_6t
Xbit_r48_c179 bl_179 br_179 wl_48 vdd gnd cell_6t
Xbit_r49_c179 bl_179 br_179 wl_49 vdd gnd cell_6t
Xbit_r50_c179 bl_179 br_179 wl_50 vdd gnd cell_6t
Xbit_r51_c179 bl_179 br_179 wl_51 vdd gnd cell_6t
Xbit_r52_c179 bl_179 br_179 wl_52 vdd gnd cell_6t
Xbit_r53_c179 bl_179 br_179 wl_53 vdd gnd cell_6t
Xbit_r54_c179 bl_179 br_179 wl_54 vdd gnd cell_6t
Xbit_r55_c179 bl_179 br_179 wl_55 vdd gnd cell_6t
Xbit_r56_c179 bl_179 br_179 wl_56 vdd gnd cell_6t
Xbit_r57_c179 bl_179 br_179 wl_57 vdd gnd cell_6t
Xbit_r58_c179 bl_179 br_179 wl_58 vdd gnd cell_6t
Xbit_r59_c179 bl_179 br_179 wl_59 vdd gnd cell_6t
Xbit_r60_c179 bl_179 br_179 wl_60 vdd gnd cell_6t
Xbit_r61_c179 bl_179 br_179 wl_61 vdd gnd cell_6t
Xbit_r62_c179 bl_179 br_179 wl_62 vdd gnd cell_6t
Xbit_r63_c179 bl_179 br_179 wl_63 vdd gnd cell_6t
Xbit_r64_c179 bl_179 br_179 wl_64 vdd gnd cell_6t
Xbit_r65_c179 bl_179 br_179 wl_65 vdd gnd cell_6t
Xbit_r66_c179 bl_179 br_179 wl_66 vdd gnd cell_6t
Xbit_r67_c179 bl_179 br_179 wl_67 vdd gnd cell_6t
Xbit_r68_c179 bl_179 br_179 wl_68 vdd gnd cell_6t
Xbit_r69_c179 bl_179 br_179 wl_69 vdd gnd cell_6t
Xbit_r70_c179 bl_179 br_179 wl_70 vdd gnd cell_6t
Xbit_r71_c179 bl_179 br_179 wl_71 vdd gnd cell_6t
Xbit_r72_c179 bl_179 br_179 wl_72 vdd gnd cell_6t
Xbit_r73_c179 bl_179 br_179 wl_73 vdd gnd cell_6t
Xbit_r74_c179 bl_179 br_179 wl_74 vdd gnd cell_6t
Xbit_r75_c179 bl_179 br_179 wl_75 vdd gnd cell_6t
Xbit_r76_c179 bl_179 br_179 wl_76 vdd gnd cell_6t
Xbit_r77_c179 bl_179 br_179 wl_77 vdd gnd cell_6t
Xbit_r78_c179 bl_179 br_179 wl_78 vdd gnd cell_6t
Xbit_r79_c179 bl_179 br_179 wl_79 vdd gnd cell_6t
Xbit_r80_c179 bl_179 br_179 wl_80 vdd gnd cell_6t
Xbit_r81_c179 bl_179 br_179 wl_81 vdd gnd cell_6t
Xbit_r82_c179 bl_179 br_179 wl_82 vdd gnd cell_6t
Xbit_r83_c179 bl_179 br_179 wl_83 vdd gnd cell_6t
Xbit_r84_c179 bl_179 br_179 wl_84 vdd gnd cell_6t
Xbit_r85_c179 bl_179 br_179 wl_85 vdd gnd cell_6t
Xbit_r86_c179 bl_179 br_179 wl_86 vdd gnd cell_6t
Xbit_r87_c179 bl_179 br_179 wl_87 vdd gnd cell_6t
Xbit_r88_c179 bl_179 br_179 wl_88 vdd gnd cell_6t
Xbit_r89_c179 bl_179 br_179 wl_89 vdd gnd cell_6t
Xbit_r90_c179 bl_179 br_179 wl_90 vdd gnd cell_6t
Xbit_r91_c179 bl_179 br_179 wl_91 vdd gnd cell_6t
Xbit_r92_c179 bl_179 br_179 wl_92 vdd gnd cell_6t
Xbit_r93_c179 bl_179 br_179 wl_93 vdd gnd cell_6t
Xbit_r94_c179 bl_179 br_179 wl_94 vdd gnd cell_6t
Xbit_r95_c179 bl_179 br_179 wl_95 vdd gnd cell_6t
Xbit_r96_c179 bl_179 br_179 wl_96 vdd gnd cell_6t
Xbit_r97_c179 bl_179 br_179 wl_97 vdd gnd cell_6t
Xbit_r98_c179 bl_179 br_179 wl_98 vdd gnd cell_6t
Xbit_r99_c179 bl_179 br_179 wl_99 vdd gnd cell_6t
Xbit_r100_c179 bl_179 br_179 wl_100 vdd gnd cell_6t
Xbit_r101_c179 bl_179 br_179 wl_101 vdd gnd cell_6t
Xbit_r102_c179 bl_179 br_179 wl_102 vdd gnd cell_6t
Xbit_r103_c179 bl_179 br_179 wl_103 vdd gnd cell_6t
Xbit_r104_c179 bl_179 br_179 wl_104 vdd gnd cell_6t
Xbit_r105_c179 bl_179 br_179 wl_105 vdd gnd cell_6t
Xbit_r106_c179 bl_179 br_179 wl_106 vdd gnd cell_6t
Xbit_r107_c179 bl_179 br_179 wl_107 vdd gnd cell_6t
Xbit_r108_c179 bl_179 br_179 wl_108 vdd gnd cell_6t
Xbit_r109_c179 bl_179 br_179 wl_109 vdd gnd cell_6t
Xbit_r110_c179 bl_179 br_179 wl_110 vdd gnd cell_6t
Xbit_r111_c179 bl_179 br_179 wl_111 vdd gnd cell_6t
Xbit_r112_c179 bl_179 br_179 wl_112 vdd gnd cell_6t
Xbit_r113_c179 bl_179 br_179 wl_113 vdd gnd cell_6t
Xbit_r114_c179 bl_179 br_179 wl_114 vdd gnd cell_6t
Xbit_r115_c179 bl_179 br_179 wl_115 vdd gnd cell_6t
Xbit_r116_c179 bl_179 br_179 wl_116 vdd gnd cell_6t
Xbit_r117_c179 bl_179 br_179 wl_117 vdd gnd cell_6t
Xbit_r118_c179 bl_179 br_179 wl_118 vdd gnd cell_6t
Xbit_r119_c179 bl_179 br_179 wl_119 vdd gnd cell_6t
Xbit_r120_c179 bl_179 br_179 wl_120 vdd gnd cell_6t
Xbit_r121_c179 bl_179 br_179 wl_121 vdd gnd cell_6t
Xbit_r122_c179 bl_179 br_179 wl_122 vdd gnd cell_6t
Xbit_r123_c179 bl_179 br_179 wl_123 vdd gnd cell_6t
Xbit_r124_c179 bl_179 br_179 wl_124 vdd gnd cell_6t
Xbit_r125_c179 bl_179 br_179 wl_125 vdd gnd cell_6t
Xbit_r126_c179 bl_179 br_179 wl_126 vdd gnd cell_6t
Xbit_r127_c179 bl_179 br_179 wl_127 vdd gnd cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd cell_6t
Xbit_r1_c180 bl_180 br_180 wl_1 vdd gnd cell_6t
Xbit_r2_c180 bl_180 br_180 wl_2 vdd gnd cell_6t
Xbit_r3_c180 bl_180 br_180 wl_3 vdd gnd cell_6t
Xbit_r4_c180 bl_180 br_180 wl_4 vdd gnd cell_6t
Xbit_r5_c180 bl_180 br_180 wl_5 vdd gnd cell_6t
Xbit_r6_c180 bl_180 br_180 wl_6 vdd gnd cell_6t
Xbit_r7_c180 bl_180 br_180 wl_7 vdd gnd cell_6t
Xbit_r8_c180 bl_180 br_180 wl_8 vdd gnd cell_6t
Xbit_r9_c180 bl_180 br_180 wl_9 vdd gnd cell_6t
Xbit_r10_c180 bl_180 br_180 wl_10 vdd gnd cell_6t
Xbit_r11_c180 bl_180 br_180 wl_11 vdd gnd cell_6t
Xbit_r12_c180 bl_180 br_180 wl_12 vdd gnd cell_6t
Xbit_r13_c180 bl_180 br_180 wl_13 vdd gnd cell_6t
Xbit_r14_c180 bl_180 br_180 wl_14 vdd gnd cell_6t
Xbit_r15_c180 bl_180 br_180 wl_15 vdd gnd cell_6t
Xbit_r16_c180 bl_180 br_180 wl_16 vdd gnd cell_6t
Xbit_r17_c180 bl_180 br_180 wl_17 vdd gnd cell_6t
Xbit_r18_c180 bl_180 br_180 wl_18 vdd gnd cell_6t
Xbit_r19_c180 bl_180 br_180 wl_19 vdd gnd cell_6t
Xbit_r20_c180 bl_180 br_180 wl_20 vdd gnd cell_6t
Xbit_r21_c180 bl_180 br_180 wl_21 vdd gnd cell_6t
Xbit_r22_c180 bl_180 br_180 wl_22 vdd gnd cell_6t
Xbit_r23_c180 bl_180 br_180 wl_23 vdd gnd cell_6t
Xbit_r24_c180 bl_180 br_180 wl_24 vdd gnd cell_6t
Xbit_r25_c180 bl_180 br_180 wl_25 vdd gnd cell_6t
Xbit_r26_c180 bl_180 br_180 wl_26 vdd gnd cell_6t
Xbit_r27_c180 bl_180 br_180 wl_27 vdd gnd cell_6t
Xbit_r28_c180 bl_180 br_180 wl_28 vdd gnd cell_6t
Xbit_r29_c180 bl_180 br_180 wl_29 vdd gnd cell_6t
Xbit_r30_c180 bl_180 br_180 wl_30 vdd gnd cell_6t
Xbit_r31_c180 bl_180 br_180 wl_31 vdd gnd cell_6t
Xbit_r32_c180 bl_180 br_180 wl_32 vdd gnd cell_6t
Xbit_r33_c180 bl_180 br_180 wl_33 vdd gnd cell_6t
Xbit_r34_c180 bl_180 br_180 wl_34 vdd gnd cell_6t
Xbit_r35_c180 bl_180 br_180 wl_35 vdd gnd cell_6t
Xbit_r36_c180 bl_180 br_180 wl_36 vdd gnd cell_6t
Xbit_r37_c180 bl_180 br_180 wl_37 vdd gnd cell_6t
Xbit_r38_c180 bl_180 br_180 wl_38 vdd gnd cell_6t
Xbit_r39_c180 bl_180 br_180 wl_39 vdd gnd cell_6t
Xbit_r40_c180 bl_180 br_180 wl_40 vdd gnd cell_6t
Xbit_r41_c180 bl_180 br_180 wl_41 vdd gnd cell_6t
Xbit_r42_c180 bl_180 br_180 wl_42 vdd gnd cell_6t
Xbit_r43_c180 bl_180 br_180 wl_43 vdd gnd cell_6t
Xbit_r44_c180 bl_180 br_180 wl_44 vdd gnd cell_6t
Xbit_r45_c180 bl_180 br_180 wl_45 vdd gnd cell_6t
Xbit_r46_c180 bl_180 br_180 wl_46 vdd gnd cell_6t
Xbit_r47_c180 bl_180 br_180 wl_47 vdd gnd cell_6t
Xbit_r48_c180 bl_180 br_180 wl_48 vdd gnd cell_6t
Xbit_r49_c180 bl_180 br_180 wl_49 vdd gnd cell_6t
Xbit_r50_c180 bl_180 br_180 wl_50 vdd gnd cell_6t
Xbit_r51_c180 bl_180 br_180 wl_51 vdd gnd cell_6t
Xbit_r52_c180 bl_180 br_180 wl_52 vdd gnd cell_6t
Xbit_r53_c180 bl_180 br_180 wl_53 vdd gnd cell_6t
Xbit_r54_c180 bl_180 br_180 wl_54 vdd gnd cell_6t
Xbit_r55_c180 bl_180 br_180 wl_55 vdd gnd cell_6t
Xbit_r56_c180 bl_180 br_180 wl_56 vdd gnd cell_6t
Xbit_r57_c180 bl_180 br_180 wl_57 vdd gnd cell_6t
Xbit_r58_c180 bl_180 br_180 wl_58 vdd gnd cell_6t
Xbit_r59_c180 bl_180 br_180 wl_59 vdd gnd cell_6t
Xbit_r60_c180 bl_180 br_180 wl_60 vdd gnd cell_6t
Xbit_r61_c180 bl_180 br_180 wl_61 vdd gnd cell_6t
Xbit_r62_c180 bl_180 br_180 wl_62 vdd gnd cell_6t
Xbit_r63_c180 bl_180 br_180 wl_63 vdd gnd cell_6t
Xbit_r64_c180 bl_180 br_180 wl_64 vdd gnd cell_6t
Xbit_r65_c180 bl_180 br_180 wl_65 vdd gnd cell_6t
Xbit_r66_c180 bl_180 br_180 wl_66 vdd gnd cell_6t
Xbit_r67_c180 bl_180 br_180 wl_67 vdd gnd cell_6t
Xbit_r68_c180 bl_180 br_180 wl_68 vdd gnd cell_6t
Xbit_r69_c180 bl_180 br_180 wl_69 vdd gnd cell_6t
Xbit_r70_c180 bl_180 br_180 wl_70 vdd gnd cell_6t
Xbit_r71_c180 bl_180 br_180 wl_71 vdd gnd cell_6t
Xbit_r72_c180 bl_180 br_180 wl_72 vdd gnd cell_6t
Xbit_r73_c180 bl_180 br_180 wl_73 vdd gnd cell_6t
Xbit_r74_c180 bl_180 br_180 wl_74 vdd gnd cell_6t
Xbit_r75_c180 bl_180 br_180 wl_75 vdd gnd cell_6t
Xbit_r76_c180 bl_180 br_180 wl_76 vdd gnd cell_6t
Xbit_r77_c180 bl_180 br_180 wl_77 vdd gnd cell_6t
Xbit_r78_c180 bl_180 br_180 wl_78 vdd gnd cell_6t
Xbit_r79_c180 bl_180 br_180 wl_79 vdd gnd cell_6t
Xbit_r80_c180 bl_180 br_180 wl_80 vdd gnd cell_6t
Xbit_r81_c180 bl_180 br_180 wl_81 vdd gnd cell_6t
Xbit_r82_c180 bl_180 br_180 wl_82 vdd gnd cell_6t
Xbit_r83_c180 bl_180 br_180 wl_83 vdd gnd cell_6t
Xbit_r84_c180 bl_180 br_180 wl_84 vdd gnd cell_6t
Xbit_r85_c180 bl_180 br_180 wl_85 vdd gnd cell_6t
Xbit_r86_c180 bl_180 br_180 wl_86 vdd gnd cell_6t
Xbit_r87_c180 bl_180 br_180 wl_87 vdd gnd cell_6t
Xbit_r88_c180 bl_180 br_180 wl_88 vdd gnd cell_6t
Xbit_r89_c180 bl_180 br_180 wl_89 vdd gnd cell_6t
Xbit_r90_c180 bl_180 br_180 wl_90 vdd gnd cell_6t
Xbit_r91_c180 bl_180 br_180 wl_91 vdd gnd cell_6t
Xbit_r92_c180 bl_180 br_180 wl_92 vdd gnd cell_6t
Xbit_r93_c180 bl_180 br_180 wl_93 vdd gnd cell_6t
Xbit_r94_c180 bl_180 br_180 wl_94 vdd gnd cell_6t
Xbit_r95_c180 bl_180 br_180 wl_95 vdd gnd cell_6t
Xbit_r96_c180 bl_180 br_180 wl_96 vdd gnd cell_6t
Xbit_r97_c180 bl_180 br_180 wl_97 vdd gnd cell_6t
Xbit_r98_c180 bl_180 br_180 wl_98 vdd gnd cell_6t
Xbit_r99_c180 bl_180 br_180 wl_99 vdd gnd cell_6t
Xbit_r100_c180 bl_180 br_180 wl_100 vdd gnd cell_6t
Xbit_r101_c180 bl_180 br_180 wl_101 vdd gnd cell_6t
Xbit_r102_c180 bl_180 br_180 wl_102 vdd gnd cell_6t
Xbit_r103_c180 bl_180 br_180 wl_103 vdd gnd cell_6t
Xbit_r104_c180 bl_180 br_180 wl_104 vdd gnd cell_6t
Xbit_r105_c180 bl_180 br_180 wl_105 vdd gnd cell_6t
Xbit_r106_c180 bl_180 br_180 wl_106 vdd gnd cell_6t
Xbit_r107_c180 bl_180 br_180 wl_107 vdd gnd cell_6t
Xbit_r108_c180 bl_180 br_180 wl_108 vdd gnd cell_6t
Xbit_r109_c180 bl_180 br_180 wl_109 vdd gnd cell_6t
Xbit_r110_c180 bl_180 br_180 wl_110 vdd gnd cell_6t
Xbit_r111_c180 bl_180 br_180 wl_111 vdd gnd cell_6t
Xbit_r112_c180 bl_180 br_180 wl_112 vdd gnd cell_6t
Xbit_r113_c180 bl_180 br_180 wl_113 vdd gnd cell_6t
Xbit_r114_c180 bl_180 br_180 wl_114 vdd gnd cell_6t
Xbit_r115_c180 bl_180 br_180 wl_115 vdd gnd cell_6t
Xbit_r116_c180 bl_180 br_180 wl_116 vdd gnd cell_6t
Xbit_r117_c180 bl_180 br_180 wl_117 vdd gnd cell_6t
Xbit_r118_c180 bl_180 br_180 wl_118 vdd gnd cell_6t
Xbit_r119_c180 bl_180 br_180 wl_119 vdd gnd cell_6t
Xbit_r120_c180 bl_180 br_180 wl_120 vdd gnd cell_6t
Xbit_r121_c180 bl_180 br_180 wl_121 vdd gnd cell_6t
Xbit_r122_c180 bl_180 br_180 wl_122 vdd gnd cell_6t
Xbit_r123_c180 bl_180 br_180 wl_123 vdd gnd cell_6t
Xbit_r124_c180 bl_180 br_180 wl_124 vdd gnd cell_6t
Xbit_r125_c180 bl_180 br_180 wl_125 vdd gnd cell_6t
Xbit_r126_c180 bl_180 br_180 wl_126 vdd gnd cell_6t
Xbit_r127_c180 bl_180 br_180 wl_127 vdd gnd cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd cell_6t
Xbit_r1_c181 bl_181 br_181 wl_1 vdd gnd cell_6t
Xbit_r2_c181 bl_181 br_181 wl_2 vdd gnd cell_6t
Xbit_r3_c181 bl_181 br_181 wl_3 vdd gnd cell_6t
Xbit_r4_c181 bl_181 br_181 wl_4 vdd gnd cell_6t
Xbit_r5_c181 bl_181 br_181 wl_5 vdd gnd cell_6t
Xbit_r6_c181 bl_181 br_181 wl_6 vdd gnd cell_6t
Xbit_r7_c181 bl_181 br_181 wl_7 vdd gnd cell_6t
Xbit_r8_c181 bl_181 br_181 wl_8 vdd gnd cell_6t
Xbit_r9_c181 bl_181 br_181 wl_9 vdd gnd cell_6t
Xbit_r10_c181 bl_181 br_181 wl_10 vdd gnd cell_6t
Xbit_r11_c181 bl_181 br_181 wl_11 vdd gnd cell_6t
Xbit_r12_c181 bl_181 br_181 wl_12 vdd gnd cell_6t
Xbit_r13_c181 bl_181 br_181 wl_13 vdd gnd cell_6t
Xbit_r14_c181 bl_181 br_181 wl_14 vdd gnd cell_6t
Xbit_r15_c181 bl_181 br_181 wl_15 vdd gnd cell_6t
Xbit_r16_c181 bl_181 br_181 wl_16 vdd gnd cell_6t
Xbit_r17_c181 bl_181 br_181 wl_17 vdd gnd cell_6t
Xbit_r18_c181 bl_181 br_181 wl_18 vdd gnd cell_6t
Xbit_r19_c181 bl_181 br_181 wl_19 vdd gnd cell_6t
Xbit_r20_c181 bl_181 br_181 wl_20 vdd gnd cell_6t
Xbit_r21_c181 bl_181 br_181 wl_21 vdd gnd cell_6t
Xbit_r22_c181 bl_181 br_181 wl_22 vdd gnd cell_6t
Xbit_r23_c181 bl_181 br_181 wl_23 vdd gnd cell_6t
Xbit_r24_c181 bl_181 br_181 wl_24 vdd gnd cell_6t
Xbit_r25_c181 bl_181 br_181 wl_25 vdd gnd cell_6t
Xbit_r26_c181 bl_181 br_181 wl_26 vdd gnd cell_6t
Xbit_r27_c181 bl_181 br_181 wl_27 vdd gnd cell_6t
Xbit_r28_c181 bl_181 br_181 wl_28 vdd gnd cell_6t
Xbit_r29_c181 bl_181 br_181 wl_29 vdd gnd cell_6t
Xbit_r30_c181 bl_181 br_181 wl_30 vdd gnd cell_6t
Xbit_r31_c181 bl_181 br_181 wl_31 vdd gnd cell_6t
Xbit_r32_c181 bl_181 br_181 wl_32 vdd gnd cell_6t
Xbit_r33_c181 bl_181 br_181 wl_33 vdd gnd cell_6t
Xbit_r34_c181 bl_181 br_181 wl_34 vdd gnd cell_6t
Xbit_r35_c181 bl_181 br_181 wl_35 vdd gnd cell_6t
Xbit_r36_c181 bl_181 br_181 wl_36 vdd gnd cell_6t
Xbit_r37_c181 bl_181 br_181 wl_37 vdd gnd cell_6t
Xbit_r38_c181 bl_181 br_181 wl_38 vdd gnd cell_6t
Xbit_r39_c181 bl_181 br_181 wl_39 vdd gnd cell_6t
Xbit_r40_c181 bl_181 br_181 wl_40 vdd gnd cell_6t
Xbit_r41_c181 bl_181 br_181 wl_41 vdd gnd cell_6t
Xbit_r42_c181 bl_181 br_181 wl_42 vdd gnd cell_6t
Xbit_r43_c181 bl_181 br_181 wl_43 vdd gnd cell_6t
Xbit_r44_c181 bl_181 br_181 wl_44 vdd gnd cell_6t
Xbit_r45_c181 bl_181 br_181 wl_45 vdd gnd cell_6t
Xbit_r46_c181 bl_181 br_181 wl_46 vdd gnd cell_6t
Xbit_r47_c181 bl_181 br_181 wl_47 vdd gnd cell_6t
Xbit_r48_c181 bl_181 br_181 wl_48 vdd gnd cell_6t
Xbit_r49_c181 bl_181 br_181 wl_49 vdd gnd cell_6t
Xbit_r50_c181 bl_181 br_181 wl_50 vdd gnd cell_6t
Xbit_r51_c181 bl_181 br_181 wl_51 vdd gnd cell_6t
Xbit_r52_c181 bl_181 br_181 wl_52 vdd gnd cell_6t
Xbit_r53_c181 bl_181 br_181 wl_53 vdd gnd cell_6t
Xbit_r54_c181 bl_181 br_181 wl_54 vdd gnd cell_6t
Xbit_r55_c181 bl_181 br_181 wl_55 vdd gnd cell_6t
Xbit_r56_c181 bl_181 br_181 wl_56 vdd gnd cell_6t
Xbit_r57_c181 bl_181 br_181 wl_57 vdd gnd cell_6t
Xbit_r58_c181 bl_181 br_181 wl_58 vdd gnd cell_6t
Xbit_r59_c181 bl_181 br_181 wl_59 vdd gnd cell_6t
Xbit_r60_c181 bl_181 br_181 wl_60 vdd gnd cell_6t
Xbit_r61_c181 bl_181 br_181 wl_61 vdd gnd cell_6t
Xbit_r62_c181 bl_181 br_181 wl_62 vdd gnd cell_6t
Xbit_r63_c181 bl_181 br_181 wl_63 vdd gnd cell_6t
Xbit_r64_c181 bl_181 br_181 wl_64 vdd gnd cell_6t
Xbit_r65_c181 bl_181 br_181 wl_65 vdd gnd cell_6t
Xbit_r66_c181 bl_181 br_181 wl_66 vdd gnd cell_6t
Xbit_r67_c181 bl_181 br_181 wl_67 vdd gnd cell_6t
Xbit_r68_c181 bl_181 br_181 wl_68 vdd gnd cell_6t
Xbit_r69_c181 bl_181 br_181 wl_69 vdd gnd cell_6t
Xbit_r70_c181 bl_181 br_181 wl_70 vdd gnd cell_6t
Xbit_r71_c181 bl_181 br_181 wl_71 vdd gnd cell_6t
Xbit_r72_c181 bl_181 br_181 wl_72 vdd gnd cell_6t
Xbit_r73_c181 bl_181 br_181 wl_73 vdd gnd cell_6t
Xbit_r74_c181 bl_181 br_181 wl_74 vdd gnd cell_6t
Xbit_r75_c181 bl_181 br_181 wl_75 vdd gnd cell_6t
Xbit_r76_c181 bl_181 br_181 wl_76 vdd gnd cell_6t
Xbit_r77_c181 bl_181 br_181 wl_77 vdd gnd cell_6t
Xbit_r78_c181 bl_181 br_181 wl_78 vdd gnd cell_6t
Xbit_r79_c181 bl_181 br_181 wl_79 vdd gnd cell_6t
Xbit_r80_c181 bl_181 br_181 wl_80 vdd gnd cell_6t
Xbit_r81_c181 bl_181 br_181 wl_81 vdd gnd cell_6t
Xbit_r82_c181 bl_181 br_181 wl_82 vdd gnd cell_6t
Xbit_r83_c181 bl_181 br_181 wl_83 vdd gnd cell_6t
Xbit_r84_c181 bl_181 br_181 wl_84 vdd gnd cell_6t
Xbit_r85_c181 bl_181 br_181 wl_85 vdd gnd cell_6t
Xbit_r86_c181 bl_181 br_181 wl_86 vdd gnd cell_6t
Xbit_r87_c181 bl_181 br_181 wl_87 vdd gnd cell_6t
Xbit_r88_c181 bl_181 br_181 wl_88 vdd gnd cell_6t
Xbit_r89_c181 bl_181 br_181 wl_89 vdd gnd cell_6t
Xbit_r90_c181 bl_181 br_181 wl_90 vdd gnd cell_6t
Xbit_r91_c181 bl_181 br_181 wl_91 vdd gnd cell_6t
Xbit_r92_c181 bl_181 br_181 wl_92 vdd gnd cell_6t
Xbit_r93_c181 bl_181 br_181 wl_93 vdd gnd cell_6t
Xbit_r94_c181 bl_181 br_181 wl_94 vdd gnd cell_6t
Xbit_r95_c181 bl_181 br_181 wl_95 vdd gnd cell_6t
Xbit_r96_c181 bl_181 br_181 wl_96 vdd gnd cell_6t
Xbit_r97_c181 bl_181 br_181 wl_97 vdd gnd cell_6t
Xbit_r98_c181 bl_181 br_181 wl_98 vdd gnd cell_6t
Xbit_r99_c181 bl_181 br_181 wl_99 vdd gnd cell_6t
Xbit_r100_c181 bl_181 br_181 wl_100 vdd gnd cell_6t
Xbit_r101_c181 bl_181 br_181 wl_101 vdd gnd cell_6t
Xbit_r102_c181 bl_181 br_181 wl_102 vdd gnd cell_6t
Xbit_r103_c181 bl_181 br_181 wl_103 vdd gnd cell_6t
Xbit_r104_c181 bl_181 br_181 wl_104 vdd gnd cell_6t
Xbit_r105_c181 bl_181 br_181 wl_105 vdd gnd cell_6t
Xbit_r106_c181 bl_181 br_181 wl_106 vdd gnd cell_6t
Xbit_r107_c181 bl_181 br_181 wl_107 vdd gnd cell_6t
Xbit_r108_c181 bl_181 br_181 wl_108 vdd gnd cell_6t
Xbit_r109_c181 bl_181 br_181 wl_109 vdd gnd cell_6t
Xbit_r110_c181 bl_181 br_181 wl_110 vdd gnd cell_6t
Xbit_r111_c181 bl_181 br_181 wl_111 vdd gnd cell_6t
Xbit_r112_c181 bl_181 br_181 wl_112 vdd gnd cell_6t
Xbit_r113_c181 bl_181 br_181 wl_113 vdd gnd cell_6t
Xbit_r114_c181 bl_181 br_181 wl_114 vdd gnd cell_6t
Xbit_r115_c181 bl_181 br_181 wl_115 vdd gnd cell_6t
Xbit_r116_c181 bl_181 br_181 wl_116 vdd gnd cell_6t
Xbit_r117_c181 bl_181 br_181 wl_117 vdd gnd cell_6t
Xbit_r118_c181 bl_181 br_181 wl_118 vdd gnd cell_6t
Xbit_r119_c181 bl_181 br_181 wl_119 vdd gnd cell_6t
Xbit_r120_c181 bl_181 br_181 wl_120 vdd gnd cell_6t
Xbit_r121_c181 bl_181 br_181 wl_121 vdd gnd cell_6t
Xbit_r122_c181 bl_181 br_181 wl_122 vdd gnd cell_6t
Xbit_r123_c181 bl_181 br_181 wl_123 vdd gnd cell_6t
Xbit_r124_c181 bl_181 br_181 wl_124 vdd gnd cell_6t
Xbit_r125_c181 bl_181 br_181 wl_125 vdd gnd cell_6t
Xbit_r126_c181 bl_181 br_181 wl_126 vdd gnd cell_6t
Xbit_r127_c181 bl_181 br_181 wl_127 vdd gnd cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd cell_6t
Xbit_r1_c182 bl_182 br_182 wl_1 vdd gnd cell_6t
Xbit_r2_c182 bl_182 br_182 wl_2 vdd gnd cell_6t
Xbit_r3_c182 bl_182 br_182 wl_3 vdd gnd cell_6t
Xbit_r4_c182 bl_182 br_182 wl_4 vdd gnd cell_6t
Xbit_r5_c182 bl_182 br_182 wl_5 vdd gnd cell_6t
Xbit_r6_c182 bl_182 br_182 wl_6 vdd gnd cell_6t
Xbit_r7_c182 bl_182 br_182 wl_7 vdd gnd cell_6t
Xbit_r8_c182 bl_182 br_182 wl_8 vdd gnd cell_6t
Xbit_r9_c182 bl_182 br_182 wl_9 vdd gnd cell_6t
Xbit_r10_c182 bl_182 br_182 wl_10 vdd gnd cell_6t
Xbit_r11_c182 bl_182 br_182 wl_11 vdd gnd cell_6t
Xbit_r12_c182 bl_182 br_182 wl_12 vdd gnd cell_6t
Xbit_r13_c182 bl_182 br_182 wl_13 vdd gnd cell_6t
Xbit_r14_c182 bl_182 br_182 wl_14 vdd gnd cell_6t
Xbit_r15_c182 bl_182 br_182 wl_15 vdd gnd cell_6t
Xbit_r16_c182 bl_182 br_182 wl_16 vdd gnd cell_6t
Xbit_r17_c182 bl_182 br_182 wl_17 vdd gnd cell_6t
Xbit_r18_c182 bl_182 br_182 wl_18 vdd gnd cell_6t
Xbit_r19_c182 bl_182 br_182 wl_19 vdd gnd cell_6t
Xbit_r20_c182 bl_182 br_182 wl_20 vdd gnd cell_6t
Xbit_r21_c182 bl_182 br_182 wl_21 vdd gnd cell_6t
Xbit_r22_c182 bl_182 br_182 wl_22 vdd gnd cell_6t
Xbit_r23_c182 bl_182 br_182 wl_23 vdd gnd cell_6t
Xbit_r24_c182 bl_182 br_182 wl_24 vdd gnd cell_6t
Xbit_r25_c182 bl_182 br_182 wl_25 vdd gnd cell_6t
Xbit_r26_c182 bl_182 br_182 wl_26 vdd gnd cell_6t
Xbit_r27_c182 bl_182 br_182 wl_27 vdd gnd cell_6t
Xbit_r28_c182 bl_182 br_182 wl_28 vdd gnd cell_6t
Xbit_r29_c182 bl_182 br_182 wl_29 vdd gnd cell_6t
Xbit_r30_c182 bl_182 br_182 wl_30 vdd gnd cell_6t
Xbit_r31_c182 bl_182 br_182 wl_31 vdd gnd cell_6t
Xbit_r32_c182 bl_182 br_182 wl_32 vdd gnd cell_6t
Xbit_r33_c182 bl_182 br_182 wl_33 vdd gnd cell_6t
Xbit_r34_c182 bl_182 br_182 wl_34 vdd gnd cell_6t
Xbit_r35_c182 bl_182 br_182 wl_35 vdd gnd cell_6t
Xbit_r36_c182 bl_182 br_182 wl_36 vdd gnd cell_6t
Xbit_r37_c182 bl_182 br_182 wl_37 vdd gnd cell_6t
Xbit_r38_c182 bl_182 br_182 wl_38 vdd gnd cell_6t
Xbit_r39_c182 bl_182 br_182 wl_39 vdd gnd cell_6t
Xbit_r40_c182 bl_182 br_182 wl_40 vdd gnd cell_6t
Xbit_r41_c182 bl_182 br_182 wl_41 vdd gnd cell_6t
Xbit_r42_c182 bl_182 br_182 wl_42 vdd gnd cell_6t
Xbit_r43_c182 bl_182 br_182 wl_43 vdd gnd cell_6t
Xbit_r44_c182 bl_182 br_182 wl_44 vdd gnd cell_6t
Xbit_r45_c182 bl_182 br_182 wl_45 vdd gnd cell_6t
Xbit_r46_c182 bl_182 br_182 wl_46 vdd gnd cell_6t
Xbit_r47_c182 bl_182 br_182 wl_47 vdd gnd cell_6t
Xbit_r48_c182 bl_182 br_182 wl_48 vdd gnd cell_6t
Xbit_r49_c182 bl_182 br_182 wl_49 vdd gnd cell_6t
Xbit_r50_c182 bl_182 br_182 wl_50 vdd gnd cell_6t
Xbit_r51_c182 bl_182 br_182 wl_51 vdd gnd cell_6t
Xbit_r52_c182 bl_182 br_182 wl_52 vdd gnd cell_6t
Xbit_r53_c182 bl_182 br_182 wl_53 vdd gnd cell_6t
Xbit_r54_c182 bl_182 br_182 wl_54 vdd gnd cell_6t
Xbit_r55_c182 bl_182 br_182 wl_55 vdd gnd cell_6t
Xbit_r56_c182 bl_182 br_182 wl_56 vdd gnd cell_6t
Xbit_r57_c182 bl_182 br_182 wl_57 vdd gnd cell_6t
Xbit_r58_c182 bl_182 br_182 wl_58 vdd gnd cell_6t
Xbit_r59_c182 bl_182 br_182 wl_59 vdd gnd cell_6t
Xbit_r60_c182 bl_182 br_182 wl_60 vdd gnd cell_6t
Xbit_r61_c182 bl_182 br_182 wl_61 vdd gnd cell_6t
Xbit_r62_c182 bl_182 br_182 wl_62 vdd gnd cell_6t
Xbit_r63_c182 bl_182 br_182 wl_63 vdd gnd cell_6t
Xbit_r64_c182 bl_182 br_182 wl_64 vdd gnd cell_6t
Xbit_r65_c182 bl_182 br_182 wl_65 vdd gnd cell_6t
Xbit_r66_c182 bl_182 br_182 wl_66 vdd gnd cell_6t
Xbit_r67_c182 bl_182 br_182 wl_67 vdd gnd cell_6t
Xbit_r68_c182 bl_182 br_182 wl_68 vdd gnd cell_6t
Xbit_r69_c182 bl_182 br_182 wl_69 vdd gnd cell_6t
Xbit_r70_c182 bl_182 br_182 wl_70 vdd gnd cell_6t
Xbit_r71_c182 bl_182 br_182 wl_71 vdd gnd cell_6t
Xbit_r72_c182 bl_182 br_182 wl_72 vdd gnd cell_6t
Xbit_r73_c182 bl_182 br_182 wl_73 vdd gnd cell_6t
Xbit_r74_c182 bl_182 br_182 wl_74 vdd gnd cell_6t
Xbit_r75_c182 bl_182 br_182 wl_75 vdd gnd cell_6t
Xbit_r76_c182 bl_182 br_182 wl_76 vdd gnd cell_6t
Xbit_r77_c182 bl_182 br_182 wl_77 vdd gnd cell_6t
Xbit_r78_c182 bl_182 br_182 wl_78 vdd gnd cell_6t
Xbit_r79_c182 bl_182 br_182 wl_79 vdd gnd cell_6t
Xbit_r80_c182 bl_182 br_182 wl_80 vdd gnd cell_6t
Xbit_r81_c182 bl_182 br_182 wl_81 vdd gnd cell_6t
Xbit_r82_c182 bl_182 br_182 wl_82 vdd gnd cell_6t
Xbit_r83_c182 bl_182 br_182 wl_83 vdd gnd cell_6t
Xbit_r84_c182 bl_182 br_182 wl_84 vdd gnd cell_6t
Xbit_r85_c182 bl_182 br_182 wl_85 vdd gnd cell_6t
Xbit_r86_c182 bl_182 br_182 wl_86 vdd gnd cell_6t
Xbit_r87_c182 bl_182 br_182 wl_87 vdd gnd cell_6t
Xbit_r88_c182 bl_182 br_182 wl_88 vdd gnd cell_6t
Xbit_r89_c182 bl_182 br_182 wl_89 vdd gnd cell_6t
Xbit_r90_c182 bl_182 br_182 wl_90 vdd gnd cell_6t
Xbit_r91_c182 bl_182 br_182 wl_91 vdd gnd cell_6t
Xbit_r92_c182 bl_182 br_182 wl_92 vdd gnd cell_6t
Xbit_r93_c182 bl_182 br_182 wl_93 vdd gnd cell_6t
Xbit_r94_c182 bl_182 br_182 wl_94 vdd gnd cell_6t
Xbit_r95_c182 bl_182 br_182 wl_95 vdd gnd cell_6t
Xbit_r96_c182 bl_182 br_182 wl_96 vdd gnd cell_6t
Xbit_r97_c182 bl_182 br_182 wl_97 vdd gnd cell_6t
Xbit_r98_c182 bl_182 br_182 wl_98 vdd gnd cell_6t
Xbit_r99_c182 bl_182 br_182 wl_99 vdd gnd cell_6t
Xbit_r100_c182 bl_182 br_182 wl_100 vdd gnd cell_6t
Xbit_r101_c182 bl_182 br_182 wl_101 vdd gnd cell_6t
Xbit_r102_c182 bl_182 br_182 wl_102 vdd gnd cell_6t
Xbit_r103_c182 bl_182 br_182 wl_103 vdd gnd cell_6t
Xbit_r104_c182 bl_182 br_182 wl_104 vdd gnd cell_6t
Xbit_r105_c182 bl_182 br_182 wl_105 vdd gnd cell_6t
Xbit_r106_c182 bl_182 br_182 wl_106 vdd gnd cell_6t
Xbit_r107_c182 bl_182 br_182 wl_107 vdd gnd cell_6t
Xbit_r108_c182 bl_182 br_182 wl_108 vdd gnd cell_6t
Xbit_r109_c182 bl_182 br_182 wl_109 vdd gnd cell_6t
Xbit_r110_c182 bl_182 br_182 wl_110 vdd gnd cell_6t
Xbit_r111_c182 bl_182 br_182 wl_111 vdd gnd cell_6t
Xbit_r112_c182 bl_182 br_182 wl_112 vdd gnd cell_6t
Xbit_r113_c182 bl_182 br_182 wl_113 vdd gnd cell_6t
Xbit_r114_c182 bl_182 br_182 wl_114 vdd gnd cell_6t
Xbit_r115_c182 bl_182 br_182 wl_115 vdd gnd cell_6t
Xbit_r116_c182 bl_182 br_182 wl_116 vdd gnd cell_6t
Xbit_r117_c182 bl_182 br_182 wl_117 vdd gnd cell_6t
Xbit_r118_c182 bl_182 br_182 wl_118 vdd gnd cell_6t
Xbit_r119_c182 bl_182 br_182 wl_119 vdd gnd cell_6t
Xbit_r120_c182 bl_182 br_182 wl_120 vdd gnd cell_6t
Xbit_r121_c182 bl_182 br_182 wl_121 vdd gnd cell_6t
Xbit_r122_c182 bl_182 br_182 wl_122 vdd gnd cell_6t
Xbit_r123_c182 bl_182 br_182 wl_123 vdd gnd cell_6t
Xbit_r124_c182 bl_182 br_182 wl_124 vdd gnd cell_6t
Xbit_r125_c182 bl_182 br_182 wl_125 vdd gnd cell_6t
Xbit_r126_c182 bl_182 br_182 wl_126 vdd gnd cell_6t
Xbit_r127_c182 bl_182 br_182 wl_127 vdd gnd cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd cell_6t
Xbit_r1_c183 bl_183 br_183 wl_1 vdd gnd cell_6t
Xbit_r2_c183 bl_183 br_183 wl_2 vdd gnd cell_6t
Xbit_r3_c183 bl_183 br_183 wl_3 vdd gnd cell_6t
Xbit_r4_c183 bl_183 br_183 wl_4 vdd gnd cell_6t
Xbit_r5_c183 bl_183 br_183 wl_5 vdd gnd cell_6t
Xbit_r6_c183 bl_183 br_183 wl_6 vdd gnd cell_6t
Xbit_r7_c183 bl_183 br_183 wl_7 vdd gnd cell_6t
Xbit_r8_c183 bl_183 br_183 wl_8 vdd gnd cell_6t
Xbit_r9_c183 bl_183 br_183 wl_9 vdd gnd cell_6t
Xbit_r10_c183 bl_183 br_183 wl_10 vdd gnd cell_6t
Xbit_r11_c183 bl_183 br_183 wl_11 vdd gnd cell_6t
Xbit_r12_c183 bl_183 br_183 wl_12 vdd gnd cell_6t
Xbit_r13_c183 bl_183 br_183 wl_13 vdd gnd cell_6t
Xbit_r14_c183 bl_183 br_183 wl_14 vdd gnd cell_6t
Xbit_r15_c183 bl_183 br_183 wl_15 vdd gnd cell_6t
Xbit_r16_c183 bl_183 br_183 wl_16 vdd gnd cell_6t
Xbit_r17_c183 bl_183 br_183 wl_17 vdd gnd cell_6t
Xbit_r18_c183 bl_183 br_183 wl_18 vdd gnd cell_6t
Xbit_r19_c183 bl_183 br_183 wl_19 vdd gnd cell_6t
Xbit_r20_c183 bl_183 br_183 wl_20 vdd gnd cell_6t
Xbit_r21_c183 bl_183 br_183 wl_21 vdd gnd cell_6t
Xbit_r22_c183 bl_183 br_183 wl_22 vdd gnd cell_6t
Xbit_r23_c183 bl_183 br_183 wl_23 vdd gnd cell_6t
Xbit_r24_c183 bl_183 br_183 wl_24 vdd gnd cell_6t
Xbit_r25_c183 bl_183 br_183 wl_25 vdd gnd cell_6t
Xbit_r26_c183 bl_183 br_183 wl_26 vdd gnd cell_6t
Xbit_r27_c183 bl_183 br_183 wl_27 vdd gnd cell_6t
Xbit_r28_c183 bl_183 br_183 wl_28 vdd gnd cell_6t
Xbit_r29_c183 bl_183 br_183 wl_29 vdd gnd cell_6t
Xbit_r30_c183 bl_183 br_183 wl_30 vdd gnd cell_6t
Xbit_r31_c183 bl_183 br_183 wl_31 vdd gnd cell_6t
Xbit_r32_c183 bl_183 br_183 wl_32 vdd gnd cell_6t
Xbit_r33_c183 bl_183 br_183 wl_33 vdd gnd cell_6t
Xbit_r34_c183 bl_183 br_183 wl_34 vdd gnd cell_6t
Xbit_r35_c183 bl_183 br_183 wl_35 vdd gnd cell_6t
Xbit_r36_c183 bl_183 br_183 wl_36 vdd gnd cell_6t
Xbit_r37_c183 bl_183 br_183 wl_37 vdd gnd cell_6t
Xbit_r38_c183 bl_183 br_183 wl_38 vdd gnd cell_6t
Xbit_r39_c183 bl_183 br_183 wl_39 vdd gnd cell_6t
Xbit_r40_c183 bl_183 br_183 wl_40 vdd gnd cell_6t
Xbit_r41_c183 bl_183 br_183 wl_41 vdd gnd cell_6t
Xbit_r42_c183 bl_183 br_183 wl_42 vdd gnd cell_6t
Xbit_r43_c183 bl_183 br_183 wl_43 vdd gnd cell_6t
Xbit_r44_c183 bl_183 br_183 wl_44 vdd gnd cell_6t
Xbit_r45_c183 bl_183 br_183 wl_45 vdd gnd cell_6t
Xbit_r46_c183 bl_183 br_183 wl_46 vdd gnd cell_6t
Xbit_r47_c183 bl_183 br_183 wl_47 vdd gnd cell_6t
Xbit_r48_c183 bl_183 br_183 wl_48 vdd gnd cell_6t
Xbit_r49_c183 bl_183 br_183 wl_49 vdd gnd cell_6t
Xbit_r50_c183 bl_183 br_183 wl_50 vdd gnd cell_6t
Xbit_r51_c183 bl_183 br_183 wl_51 vdd gnd cell_6t
Xbit_r52_c183 bl_183 br_183 wl_52 vdd gnd cell_6t
Xbit_r53_c183 bl_183 br_183 wl_53 vdd gnd cell_6t
Xbit_r54_c183 bl_183 br_183 wl_54 vdd gnd cell_6t
Xbit_r55_c183 bl_183 br_183 wl_55 vdd gnd cell_6t
Xbit_r56_c183 bl_183 br_183 wl_56 vdd gnd cell_6t
Xbit_r57_c183 bl_183 br_183 wl_57 vdd gnd cell_6t
Xbit_r58_c183 bl_183 br_183 wl_58 vdd gnd cell_6t
Xbit_r59_c183 bl_183 br_183 wl_59 vdd gnd cell_6t
Xbit_r60_c183 bl_183 br_183 wl_60 vdd gnd cell_6t
Xbit_r61_c183 bl_183 br_183 wl_61 vdd gnd cell_6t
Xbit_r62_c183 bl_183 br_183 wl_62 vdd gnd cell_6t
Xbit_r63_c183 bl_183 br_183 wl_63 vdd gnd cell_6t
Xbit_r64_c183 bl_183 br_183 wl_64 vdd gnd cell_6t
Xbit_r65_c183 bl_183 br_183 wl_65 vdd gnd cell_6t
Xbit_r66_c183 bl_183 br_183 wl_66 vdd gnd cell_6t
Xbit_r67_c183 bl_183 br_183 wl_67 vdd gnd cell_6t
Xbit_r68_c183 bl_183 br_183 wl_68 vdd gnd cell_6t
Xbit_r69_c183 bl_183 br_183 wl_69 vdd gnd cell_6t
Xbit_r70_c183 bl_183 br_183 wl_70 vdd gnd cell_6t
Xbit_r71_c183 bl_183 br_183 wl_71 vdd gnd cell_6t
Xbit_r72_c183 bl_183 br_183 wl_72 vdd gnd cell_6t
Xbit_r73_c183 bl_183 br_183 wl_73 vdd gnd cell_6t
Xbit_r74_c183 bl_183 br_183 wl_74 vdd gnd cell_6t
Xbit_r75_c183 bl_183 br_183 wl_75 vdd gnd cell_6t
Xbit_r76_c183 bl_183 br_183 wl_76 vdd gnd cell_6t
Xbit_r77_c183 bl_183 br_183 wl_77 vdd gnd cell_6t
Xbit_r78_c183 bl_183 br_183 wl_78 vdd gnd cell_6t
Xbit_r79_c183 bl_183 br_183 wl_79 vdd gnd cell_6t
Xbit_r80_c183 bl_183 br_183 wl_80 vdd gnd cell_6t
Xbit_r81_c183 bl_183 br_183 wl_81 vdd gnd cell_6t
Xbit_r82_c183 bl_183 br_183 wl_82 vdd gnd cell_6t
Xbit_r83_c183 bl_183 br_183 wl_83 vdd gnd cell_6t
Xbit_r84_c183 bl_183 br_183 wl_84 vdd gnd cell_6t
Xbit_r85_c183 bl_183 br_183 wl_85 vdd gnd cell_6t
Xbit_r86_c183 bl_183 br_183 wl_86 vdd gnd cell_6t
Xbit_r87_c183 bl_183 br_183 wl_87 vdd gnd cell_6t
Xbit_r88_c183 bl_183 br_183 wl_88 vdd gnd cell_6t
Xbit_r89_c183 bl_183 br_183 wl_89 vdd gnd cell_6t
Xbit_r90_c183 bl_183 br_183 wl_90 vdd gnd cell_6t
Xbit_r91_c183 bl_183 br_183 wl_91 vdd gnd cell_6t
Xbit_r92_c183 bl_183 br_183 wl_92 vdd gnd cell_6t
Xbit_r93_c183 bl_183 br_183 wl_93 vdd gnd cell_6t
Xbit_r94_c183 bl_183 br_183 wl_94 vdd gnd cell_6t
Xbit_r95_c183 bl_183 br_183 wl_95 vdd gnd cell_6t
Xbit_r96_c183 bl_183 br_183 wl_96 vdd gnd cell_6t
Xbit_r97_c183 bl_183 br_183 wl_97 vdd gnd cell_6t
Xbit_r98_c183 bl_183 br_183 wl_98 vdd gnd cell_6t
Xbit_r99_c183 bl_183 br_183 wl_99 vdd gnd cell_6t
Xbit_r100_c183 bl_183 br_183 wl_100 vdd gnd cell_6t
Xbit_r101_c183 bl_183 br_183 wl_101 vdd gnd cell_6t
Xbit_r102_c183 bl_183 br_183 wl_102 vdd gnd cell_6t
Xbit_r103_c183 bl_183 br_183 wl_103 vdd gnd cell_6t
Xbit_r104_c183 bl_183 br_183 wl_104 vdd gnd cell_6t
Xbit_r105_c183 bl_183 br_183 wl_105 vdd gnd cell_6t
Xbit_r106_c183 bl_183 br_183 wl_106 vdd gnd cell_6t
Xbit_r107_c183 bl_183 br_183 wl_107 vdd gnd cell_6t
Xbit_r108_c183 bl_183 br_183 wl_108 vdd gnd cell_6t
Xbit_r109_c183 bl_183 br_183 wl_109 vdd gnd cell_6t
Xbit_r110_c183 bl_183 br_183 wl_110 vdd gnd cell_6t
Xbit_r111_c183 bl_183 br_183 wl_111 vdd gnd cell_6t
Xbit_r112_c183 bl_183 br_183 wl_112 vdd gnd cell_6t
Xbit_r113_c183 bl_183 br_183 wl_113 vdd gnd cell_6t
Xbit_r114_c183 bl_183 br_183 wl_114 vdd gnd cell_6t
Xbit_r115_c183 bl_183 br_183 wl_115 vdd gnd cell_6t
Xbit_r116_c183 bl_183 br_183 wl_116 vdd gnd cell_6t
Xbit_r117_c183 bl_183 br_183 wl_117 vdd gnd cell_6t
Xbit_r118_c183 bl_183 br_183 wl_118 vdd gnd cell_6t
Xbit_r119_c183 bl_183 br_183 wl_119 vdd gnd cell_6t
Xbit_r120_c183 bl_183 br_183 wl_120 vdd gnd cell_6t
Xbit_r121_c183 bl_183 br_183 wl_121 vdd gnd cell_6t
Xbit_r122_c183 bl_183 br_183 wl_122 vdd gnd cell_6t
Xbit_r123_c183 bl_183 br_183 wl_123 vdd gnd cell_6t
Xbit_r124_c183 bl_183 br_183 wl_124 vdd gnd cell_6t
Xbit_r125_c183 bl_183 br_183 wl_125 vdd gnd cell_6t
Xbit_r126_c183 bl_183 br_183 wl_126 vdd gnd cell_6t
Xbit_r127_c183 bl_183 br_183 wl_127 vdd gnd cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd cell_6t
Xbit_r1_c184 bl_184 br_184 wl_1 vdd gnd cell_6t
Xbit_r2_c184 bl_184 br_184 wl_2 vdd gnd cell_6t
Xbit_r3_c184 bl_184 br_184 wl_3 vdd gnd cell_6t
Xbit_r4_c184 bl_184 br_184 wl_4 vdd gnd cell_6t
Xbit_r5_c184 bl_184 br_184 wl_5 vdd gnd cell_6t
Xbit_r6_c184 bl_184 br_184 wl_6 vdd gnd cell_6t
Xbit_r7_c184 bl_184 br_184 wl_7 vdd gnd cell_6t
Xbit_r8_c184 bl_184 br_184 wl_8 vdd gnd cell_6t
Xbit_r9_c184 bl_184 br_184 wl_9 vdd gnd cell_6t
Xbit_r10_c184 bl_184 br_184 wl_10 vdd gnd cell_6t
Xbit_r11_c184 bl_184 br_184 wl_11 vdd gnd cell_6t
Xbit_r12_c184 bl_184 br_184 wl_12 vdd gnd cell_6t
Xbit_r13_c184 bl_184 br_184 wl_13 vdd gnd cell_6t
Xbit_r14_c184 bl_184 br_184 wl_14 vdd gnd cell_6t
Xbit_r15_c184 bl_184 br_184 wl_15 vdd gnd cell_6t
Xbit_r16_c184 bl_184 br_184 wl_16 vdd gnd cell_6t
Xbit_r17_c184 bl_184 br_184 wl_17 vdd gnd cell_6t
Xbit_r18_c184 bl_184 br_184 wl_18 vdd gnd cell_6t
Xbit_r19_c184 bl_184 br_184 wl_19 vdd gnd cell_6t
Xbit_r20_c184 bl_184 br_184 wl_20 vdd gnd cell_6t
Xbit_r21_c184 bl_184 br_184 wl_21 vdd gnd cell_6t
Xbit_r22_c184 bl_184 br_184 wl_22 vdd gnd cell_6t
Xbit_r23_c184 bl_184 br_184 wl_23 vdd gnd cell_6t
Xbit_r24_c184 bl_184 br_184 wl_24 vdd gnd cell_6t
Xbit_r25_c184 bl_184 br_184 wl_25 vdd gnd cell_6t
Xbit_r26_c184 bl_184 br_184 wl_26 vdd gnd cell_6t
Xbit_r27_c184 bl_184 br_184 wl_27 vdd gnd cell_6t
Xbit_r28_c184 bl_184 br_184 wl_28 vdd gnd cell_6t
Xbit_r29_c184 bl_184 br_184 wl_29 vdd gnd cell_6t
Xbit_r30_c184 bl_184 br_184 wl_30 vdd gnd cell_6t
Xbit_r31_c184 bl_184 br_184 wl_31 vdd gnd cell_6t
Xbit_r32_c184 bl_184 br_184 wl_32 vdd gnd cell_6t
Xbit_r33_c184 bl_184 br_184 wl_33 vdd gnd cell_6t
Xbit_r34_c184 bl_184 br_184 wl_34 vdd gnd cell_6t
Xbit_r35_c184 bl_184 br_184 wl_35 vdd gnd cell_6t
Xbit_r36_c184 bl_184 br_184 wl_36 vdd gnd cell_6t
Xbit_r37_c184 bl_184 br_184 wl_37 vdd gnd cell_6t
Xbit_r38_c184 bl_184 br_184 wl_38 vdd gnd cell_6t
Xbit_r39_c184 bl_184 br_184 wl_39 vdd gnd cell_6t
Xbit_r40_c184 bl_184 br_184 wl_40 vdd gnd cell_6t
Xbit_r41_c184 bl_184 br_184 wl_41 vdd gnd cell_6t
Xbit_r42_c184 bl_184 br_184 wl_42 vdd gnd cell_6t
Xbit_r43_c184 bl_184 br_184 wl_43 vdd gnd cell_6t
Xbit_r44_c184 bl_184 br_184 wl_44 vdd gnd cell_6t
Xbit_r45_c184 bl_184 br_184 wl_45 vdd gnd cell_6t
Xbit_r46_c184 bl_184 br_184 wl_46 vdd gnd cell_6t
Xbit_r47_c184 bl_184 br_184 wl_47 vdd gnd cell_6t
Xbit_r48_c184 bl_184 br_184 wl_48 vdd gnd cell_6t
Xbit_r49_c184 bl_184 br_184 wl_49 vdd gnd cell_6t
Xbit_r50_c184 bl_184 br_184 wl_50 vdd gnd cell_6t
Xbit_r51_c184 bl_184 br_184 wl_51 vdd gnd cell_6t
Xbit_r52_c184 bl_184 br_184 wl_52 vdd gnd cell_6t
Xbit_r53_c184 bl_184 br_184 wl_53 vdd gnd cell_6t
Xbit_r54_c184 bl_184 br_184 wl_54 vdd gnd cell_6t
Xbit_r55_c184 bl_184 br_184 wl_55 vdd gnd cell_6t
Xbit_r56_c184 bl_184 br_184 wl_56 vdd gnd cell_6t
Xbit_r57_c184 bl_184 br_184 wl_57 vdd gnd cell_6t
Xbit_r58_c184 bl_184 br_184 wl_58 vdd gnd cell_6t
Xbit_r59_c184 bl_184 br_184 wl_59 vdd gnd cell_6t
Xbit_r60_c184 bl_184 br_184 wl_60 vdd gnd cell_6t
Xbit_r61_c184 bl_184 br_184 wl_61 vdd gnd cell_6t
Xbit_r62_c184 bl_184 br_184 wl_62 vdd gnd cell_6t
Xbit_r63_c184 bl_184 br_184 wl_63 vdd gnd cell_6t
Xbit_r64_c184 bl_184 br_184 wl_64 vdd gnd cell_6t
Xbit_r65_c184 bl_184 br_184 wl_65 vdd gnd cell_6t
Xbit_r66_c184 bl_184 br_184 wl_66 vdd gnd cell_6t
Xbit_r67_c184 bl_184 br_184 wl_67 vdd gnd cell_6t
Xbit_r68_c184 bl_184 br_184 wl_68 vdd gnd cell_6t
Xbit_r69_c184 bl_184 br_184 wl_69 vdd gnd cell_6t
Xbit_r70_c184 bl_184 br_184 wl_70 vdd gnd cell_6t
Xbit_r71_c184 bl_184 br_184 wl_71 vdd gnd cell_6t
Xbit_r72_c184 bl_184 br_184 wl_72 vdd gnd cell_6t
Xbit_r73_c184 bl_184 br_184 wl_73 vdd gnd cell_6t
Xbit_r74_c184 bl_184 br_184 wl_74 vdd gnd cell_6t
Xbit_r75_c184 bl_184 br_184 wl_75 vdd gnd cell_6t
Xbit_r76_c184 bl_184 br_184 wl_76 vdd gnd cell_6t
Xbit_r77_c184 bl_184 br_184 wl_77 vdd gnd cell_6t
Xbit_r78_c184 bl_184 br_184 wl_78 vdd gnd cell_6t
Xbit_r79_c184 bl_184 br_184 wl_79 vdd gnd cell_6t
Xbit_r80_c184 bl_184 br_184 wl_80 vdd gnd cell_6t
Xbit_r81_c184 bl_184 br_184 wl_81 vdd gnd cell_6t
Xbit_r82_c184 bl_184 br_184 wl_82 vdd gnd cell_6t
Xbit_r83_c184 bl_184 br_184 wl_83 vdd gnd cell_6t
Xbit_r84_c184 bl_184 br_184 wl_84 vdd gnd cell_6t
Xbit_r85_c184 bl_184 br_184 wl_85 vdd gnd cell_6t
Xbit_r86_c184 bl_184 br_184 wl_86 vdd gnd cell_6t
Xbit_r87_c184 bl_184 br_184 wl_87 vdd gnd cell_6t
Xbit_r88_c184 bl_184 br_184 wl_88 vdd gnd cell_6t
Xbit_r89_c184 bl_184 br_184 wl_89 vdd gnd cell_6t
Xbit_r90_c184 bl_184 br_184 wl_90 vdd gnd cell_6t
Xbit_r91_c184 bl_184 br_184 wl_91 vdd gnd cell_6t
Xbit_r92_c184 bl_184 br_184 wl_92 vdd gnd cell_6t
Xbit_r93_c184 bl_184 br_184 wl_93 vdd gnd cell_6t
Xbit_r94_c184 bl_184 br_184 wl_94 vdd gnd cell_6t
Xbit_r95_c184 bl_184 br_184 wl_95 vdd gnd cell_6t
Xbit_r96_c184 bl_184 br_184 wl_96 vdd gnd cell_6t
Xbit_r97_c184 bl_184 br_184 wl_97 vdd gnd cell_6t
Xbit_r98_c184 bl_184 br_184 wl_98 vdd gnd cell_6t
Xbit_r99_c184 bl_184 br_184 wl_99 vdd gnd cell_6t
Xbit_r100_c184 bl_184 br_184 wl_100 vdd gnd cell_6t
Xbit_r101_c184 bl_184 br_184 wl_101 vdd gnd cell_6t
Xbit_r102_c184 bl_184 br_184 wl_102 vdd gnd cell_6t
Xbit_r103_c184 bl_184 br_184 wl_103 vdd gnd cell_6t
Xbit_r104_c184 bl_184 br_184 wl_104 vdd gnd cell_6t
Xbit_r105_c184 bl_184 br_184 wl_105 vdd gnd cell_6t
Xbit_r106_c184 bl_184 br_184 wl_106 vdd gnd cell_6t
Xbit_r107_c184 bl_184 br_184 wl_107 vdd gnd cell_6t
Xbit_r108_c184 bl_184 br_184 wl_108 vdd gnd cell_6t
Xbit_r109_c184 bl_184 br_184 wl_109 vdd gnd cell_6t
Xbit_r110_c184 bl_184 br_184 wl_110 vdd gnd cell_6t
Xbit_r111_c184 bl_184 br_184 wl_111 vdd gnd cell_6t
Xbit_r112_c184 bl_184 br_184 wl_112 vdd gnd cell_6t
Xbit_r113_c184 bl_184 br_184 wl_113 vdd gnd cell_6t
Xbit_r114_c184 bl_184 br_184 wl_114 vdd gnd cell_6t
Xbit_r115_c184 bl_184 br_184 wl_115 vdd gnd cell_6t
Xbit_r116_c184 bl_184 br_184 wl_116 vdd gnd cell_6t
Xbit_r117_c184 bl_184 br_184 wl_117 vdd gnd cell_6t
Xbit_r118_c184 bl_184 br_184 wl_118 vdd gnd cell_6t
Xbit_r119_c184 bl_184 br_184 wl_119 vdd gnd cell_6t
Xbit_r120_c184 bl_184 br_184 wl_120 vdd gnd cell_6t
Xbit_r121_c184 bl_184 br_184 wl_121 vdd gnd cell_6t
Xbit_r122_c184 bl_184 br_184 wl_122 vdd gnd cell_6t
Xbit_r123_c184 bl_184 br_184 wl_123 vdd gnd cell_6t
Xbit_r124_c184 bl_184 br_184 wl_124 vdd gnd cell_6t
Xbit_r125_c184 bl_184 br_184 wl_125 vdd gnd cell_6t
Xbit_r126_c184 bl_184 br_184 wl_126 vdd gnd cell_6t
Xbit_r127_c184 bl_184 br_184 wl_127 vdd gnd cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd cell_6t
Xbit_r1_c185 bl_185 br_185 wl_1 vdd gnd cell_6t
Xbit_r2_c185 bl_185 br_185 wl_2 vdd gnd cell_6t
Xbit_r3_c185 bl_185 br_185 wl_3 vdd gnd cell_6t
Xbit_r4_c185 bl_185 br_185 wl_4 vdd gnd cell_6t
Xbit_r5_c185 bl_185 br_185 wl_5 vdd gnd cell_6t
Xbit_r6_c185 bl_185 br_185 wl_6 vdd gnd cell_6t
Xbit_r7_c185 bl_185 br_185 wl_7 vdd gnd cell_6t
Xbit_r8_c185 bl_185 br_185 wl_8 vdd gnd cell_6t
Xbit_r9_c185 bl_185 br_185 wl_9 vdd gnd cell_6t
Xbit_r10_c185 bl_185 br_185 wl_10 vdd gnd cell_6t
Xbit_r11_c185 bl_185 br_185 wl_11 vdd gnd cell_6t
Xbit_r12_c185 bl_185 br_185 wl_12 vdd gnd cell_6t
Xbit_r13_c185 bl_185 br_185 wl_13 vdd gnd cell_6t
Xbit_r14_c185 bl_185 br_185 wl_14 vdd gnd cell_6t
Xbit_r15_c185 bl_185 br_185 wl_15 vdd gnd cell_6t
Xbit_r16_c185 bl_185 br_185 wl_16 vdd gnd cell_6t
Xbit_r17_c185 bl_185 br_185 wl_17 vdd gnd cell_6t
Xbit_r18_c185 bl_185 br_185 wl_18 vdd gnd cell_6t
Xbit_r19_c185 bl_185 br_185 wl_19 vdd gnd cell_6t
Xbit_r20_c185 bl_185 br_185 wl_20 vdd gnd cell_6t
Xbit_r21_c185 bl_185 br_185 wl_21 vdd gnd cell_6t
Xbit_r22_c185 bl_185 br_185 wl_22 vdd gnd cell_6t
Xbit_r23_c185 bl_185 br_185 wl_23 vdd gnd cell_6t
Xbit_r24_c185 bl_185 br_185 wl_24 vdd gnd cell_6t
Xbit_r25_c185 bl_185 br_185 wl_25 vdd gnd cell_6t
Xbit_r26_c185 bl_185 br_185 wl_26 vdd gnd cell_6t
Xbit_r27_c185 bl_185 br_185 wl_27 vdd gnd cell_6t
Xbit_r28_c185 bl_185 br_185 wl_28 vdd gnd cell_6t
Xbit_r29_c185 bl_185 br_185 wl_29 vdd gnd cell_6t
Xbit_r30_c185 bl_185 br_185 wl_30 vdd gnd cell_6t
Xbit_r31_c185 bl_185 br_185 wl_31 vdd gnd cell_6t
Xbit_r32_c185 bl_185 br_185 wl_32 vdd gnd cell_6t
Xbit_r33_c185 bl_185 br_185 wl_33 vdd gnd cell_6t
Xbit_r34_c185 bl_185 br_185 wl_34 vdd gnd cell_6t
Xbit_r35_c185 bl_185 br_185 wl_35 vdd gnd cell_6t
Xbit_r36_c185 bl_185 br_185 wl_36 vdd gnd cell_6t
Xbit_r37_c185 bl_185 br_185 wl_37 vdd gnd cell_6t
Xbit_r38_c185 bl_185 br_185 wl_38 vdd gnd cell_6t
Xbit_r39_c185 bl_185 br_185 wl_39 vdd gnd cell_6t
Xbit_r40_c185 bl_185 br_185 wl_40 vdd gnd cell_6t
Xbit_r41_c185 bl_185 br_185 wl_41 vdd gnd cell_6t
Xbit_r42_c185 bl_185 br_185 wl_42 vdd gnd cell_6t
Xbit_r43_c185 bl_185 br_185 wl_43 vdd gnd cell_6t
Xbit_r44_c185 bl_185 br_185 wl_44 vdd gnd cell_6t
Xbit_r45_c185 bl_185 br_185 wl_45 vdd gnd cell_6t
Xbit_r46_c185 bl_185 br_185 wl_46 vdd gnd cell_6t
Xbit_r47_c185 bl_185 br_185 wl_47 vdd gnd cell_6t
Xbit_r48_c185 bl_185 br_185 wl_48 vdd gnd cell_6t
Xbit_r49_c185 bl_185 br_185 wl_49 vdd gnd cell_6t
Xbit_r50_c185 bl_185 br_185 wl_50 vdd gnd cell_6t
Xbit_r51_c185 bl_185 br_185 wl_51 vdd gnd cell_6t
Xbit_r52_c185 bl_185 br_185 wl_52 vdd gnd cell_6t
Xbit_r53_c185 bl_185 br_185 wl_53 vdd gnd cell_6t
Xbit_r54_c185 bl_185 br_185 wl_54 vdd gnd cell_6t
Xbit_r55_c185 bl_185 br_185 wl_55 vdd gnd cell_6t
Xbit_r56_c185 bl_185 br_185 wl_56 vdd gnd cell_6t
Xbit_r57_c185 bl_185 br_185 wl_57 vdd gnd cell_6t
Xbit_r58_c185 bl_185 br_185 wl_58 vdd gnd cell_6t
Xbit_r59_c185 bl_185 br_185 wl_59 vdd gnd cell_6t
Xbit_r60_c185 bl_185 br_185 wl_60 vdd gnd cell_6t
Xbit_r61_c185 bl_185 br_185 wl_61 vdd gnd cell_6t
Xbit_r62_c185 bl_185 br_185 wl_62 vdd gnd cell_6t
Xbit_r63_c185 bl_185 br_185 wl_63 vdd gnd cell_6t
Xbit_r64_c185 bl_185 br_185 wl_64 vdd gnd cell_6t
Xbit_r65_c185 bl_185 br_185 wl_65 vdd gnd cell_6t
Xbit_r66_c185 bl_185 br_185 wl_66 vdd gnd cell_6t
Xbit_r67_c185 bl_185 br_185 wl_67 vdd gnd cell_6t
Xbit_r68_c185 bl_185 br_185 wl_68 vdd gnd cell_6t
Xbit_r69_c185 bl_185 br_185 wl_69 vdd gnd cell_6t
Xbit_r70_c185 bl_185 br_185 wl_70 vdd gnd cell_6t
Xbit_r71_c185 bl_185 br_185 wl_71 vdd gnd cell_6t
Xbit_r72_c185 bl_185 br_185 wl_72 vdd gnd cell_6t
Xbit_r73_c185 bl_185 br_185 wl_73 vdd gnd cell_6t
Xbit_r74_c185 bl_185 br_185 wl_74 vdd gnd cell_6t
Xbit_r75_c185 bl_185 br_185 wl_75 vdd gnd cell_6t
Xbit_r76_c185 bl_185 br_185 wl_76 vdd gnd cell_6t
Xbit_r77_c185 bl_185 br_185 wl_77 vdd gnd cell_6t
Xbit_r78_c185 bl_185 br_185 wl_78 vdd gnd cell_6t
Xbit_r79_c185 bl_185 br_185 wl_79 vdd gnd cell_6t
Xbit_r80_c185 bl_185 br_185 wl_80 vdd gnd cell_6t
Xbit_r81_c185 bl_185 br_185 wl_81 vdd gnd cell_6t
Xbit_r82_c185 bl_185 br_185 wl_82 vdd gnd cell_6t
Xbit_r83_c185 bl_185 br_185 wl_83 vdd gnd cell_6t
Xbit_r84_c185 bl_185 br_185 wl_84 vdd gnd cell_6t
Xbit_r85_c185 bl_185 br_185 wl_85 vdd gnd cell_6t
Xbit_r86_c185 bl_185 br_185 wl_86 vdd gnd cell_6t
Xbit_r87_c185 bl_185 br_185 wl_87 vdd gnd cell_6t
Xbit_r88_c185 bl_185 br_185 wl_88 vdd gnd cell_6t
Xbit_r89_c185 bl_185 br_185 wl_89 vdd gnd cell_6t
Xbit_r90_c185 bl_185 br_185 wl_90 vdd gnd cell_6t
Xbit_r91_c185 bl_185 br_185 wl_91 vdd gnd cell_6t
Xbit_r92_c185 bl_185 br_185 wl_92 vdd gnd cell_6t
Xbit_r93_c185 bl_185 br_185 wl_93 vdd gnd cell_6t
Xbit_r94_c185 bl_185 br_185 wl_94 vdd gnd cell_6t
Xbit_r95_c185 bl_185 br_185 wl_95 vdd gnd cell_6t
Xbit_r96_c185 bl_185 br_185 wl_96 vdd gnd cell_6t
Xbit_r97_c185 bl_185 br_185 wl_97 vdd gnd cell_6t
Xbit_r98_c185 bl_185 br_185 wl_98 vdd gnd cell_6t
Xbit_r99_c185 bl_185 br_185 wl_99 vdd gnd cell_6t
Xbit_r100_c185 bl_185 br_185 wl_100 vdd gnd cell_6t
Xbit_r101_c185 bl_185 br_185 wl_101 vdd gnd cell_6t
Xbit_r102_c185 bl_185 br_185 wl_102 vdd gnd cell_6t
Xbit_r103_c185 bl_185 br_185 wl_103 vdd gnd cell_6t
Xbit_r104_c185 bl_185 br_185 wl_104 vdd gnd cell_6t
Xbit_r105_c185 bl_185 br_185 wl_105 vdd gnd cell_6t
Xbit_r106_c185 bl_185 br_185 wl_106 vdd gnd cell_6t
Xbit_r107_c185 bl_185 br_185 wl_107 vdd gnd cell_6t
Xbit_r108_c185 bl_185 br_185 wl_108 vdd gnd cell_6t
Xbit_r109_c185 bl_185 br_185 wl_109 vdd gnd cell_6t
Xbit_r110_c185 bl_185 br_185 wl_110 vdd gnd cell_6t
Xbit_r111_c185 bl_185 br_185 wl_111 vdd gnd cell_6t
Xbit_r112_c185 bl_185 br_185 wl_112 vdd gnd cell_6t
Xbit_r113_c185 bl_185 br_185 wl_113 vdd gnd cell_6t
Xbit_r114_c185 bl_185 br_185 wl_114 vdd gnd cell_6t
Xbit_r115_c185 bl_185 br_185 wl_115 vdd gnd cell_6t
Xbit_r116_c185 bl_185 br_185 wl_116 vdd gnd cell_6t
Xbit_r117_c185 bl_185 br_185 wl_117 vdd gnd cell_6t
Xbit_r118_c185 bl_185 br_185 wl_118 vdd gnd cell_6t
Xbit_r119_c185 bl_185 br_185 wl_119 vdd gnd cell_6t
Xbit_r120_c185 bl_185 br_185 wl_120 vdd gnd cell_6t
Xbit_r121_c185 bl_185 br_185 wl_121 vdd gnd cell_6t
Xbit_r122_c185 bl_185 br_185 wl_122 vdd gnd cell_6t
Xbit_r123_c185 bl_185 br_185 wl_123 vdd gnd cell_6t
Xbit_r124_c185 bl_185 br_185 wl_124 vdd gnd cell_6t
Xbit_r125_c185 bl_185 br_185 wl_125 vdd gnd cell_6t
Xbit_r126_c185 bl_185 br_185 wl_126 vdd gnd cell_6t
Xbit_r127_c185 bl_185 br_185 wl_127 vdd gnd cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd cell_6t
Xbit_r1_c186 bl_186 br_186 wl_1 vdd gnd cell_6t
Xbit_r2_c186 bl_186 br_186 wl_2 vdd gnd cell_6t
Xbit_r3_c186 bl_186 br_186 wl_3 vdd gnd cell_6t
Xbit_r4_c186 bl_186 br_186 wl_4 vdd gnd cell_6t
Xbit_r5_c186 bl_186 br_186 wl_5 vdd gnd cell_6t
Xbit_r6_c186 bl_186 br_186 wl_6 vdd gnd cell_6t
Xbit_r7_c186 bl_186 br_186 wl_7 vdd gnd cell_6t
Xbit_r8_c186 bl_186 br_186 wl_8 vdd gnd cell_6t
Xbit_r9_c186 bl_186 br_186 wl_9 vdd gnd cell_6t
Xbit_r10_c186 bl_186 br_186 wl_10 vdd gnd cell_6t
Xbit_r11_c186 bl_186 br_186 wl_11 vdd gnd cell_6t
Xbit_r12_c186 bl_186 br_186 wl_12 vdd gnd cell_6t
Xbit_r13_c186 bl_186 br_186 wl_13 vdd gnd cell_6t
Xbit_r14_c186 bl_186 br_186 wl_14 vdd gnd cell_6t
Xbit_r15_c186 bl_186 br_186 wl_15 vdd gnd cell_6t
Xbit_r16_c186 bl_186 br_186 wl_16 vdd gnd cell_6t
Xbit_r17_c186 bl_186 br_186 wl_17 vdd gnd cell_6t
Xbit_r18_c186 bl_186 br_186 wl_18 vdd gnd cell_6t
Xbit_r19_c186 bl_186 br_186 wl_19 vdd gnd cell_6t
Xbit_r20_c186 bl_186 br_186 wl_20 vdd gnd cell_6t
Xbit_r21_c186 bl_186 br_186 wl_21 vdd gnd cell_6t
Xbit_r22_c186 bl_186 br_186 wl_22 vdd gnd cell_6t
Xbit_r23_c186 bl_186 br_186 wl_23 vdd gnd cell_6t
Xbit_r24_c186 bl_186 br_186 wl_24 vdd gnd cell_6t
Xbit_r25_c186 bl_186 br_186 wl_25 vdd gnd cell_6t
Xbit_r26_c186 bl_186 br_186 wl_26 vdd gnd cell_6t
Xbit_r27_c186 bl_186 br_186 wl_27 vdd gnd cell_6t
Xbit_r28_c186 bl_186 br_186 wl_28 vdd gnd cell_6t
Xbit_r29_c186 bl_186 br_186 wl_29 vdd gnd cell_6t
Xbit_r30_c186 bl_186 br_186 wl_30 vdd gnd cell_6t
Xbit_r31_c186 bl_186 br_186 wl_31 vdd gnd cell_6t
Xbit_r32_c186 bl_186 br_186 wl_32 vdd gnd cell_6t
Xbit_r33_c186 bl_186 br_186 wl_33 vdd gnd cell_6t
Xbit_r34_c186 bl_186 br_186 wl_34 vdd gnd cell_6t
Xbit_r35_c186 bl_186 br_186 wl_35 vdd gnd cell_6t
Xbit_r36_c186 bl_186 br_186 wl_36 vdd gnd cell_6t
Xbit_r37_c186 bl_186 br_186 wl_37 vdd gnd cell_6t
Xbit_r38_c186 bl_186 br_186 wl_38 vdd gnd cell_6t
Xbit_r39_c186 bl_186 br_186 wl_39 vdd gnd cell_6t
Xbit_r40_c186 bl_186 br_186 wl_40 vdd gnd cell_6t
Xbit_r41_c186 bl_186 br_186 wl_41 vdd gnd cell_6t
Xbit_r42_c186 bl_186 br_186 wl_42 vdd gnd cell_6t
Xbit_r43_c186 bl_186 br_186 wl_43 vdd gnd cell_6t
Xbit_r44_c186 bl_186 br_186 wl_44 vdd gnd cell_6t
Xbit_r45_c186 bl_186 br_186 wl_45 vdd gnd cell_6t
Xbit_r46_c186 bl_186 br_186 wl_46 vdd gnd cell_6t
Xbit_r47_c186 bl_186 br_186 wl_47 vdd gnd cell_6t
Xbit_r48_c186 bl_186 br_186 wl_48 vdd gnd cell_6t
Xbit_r49_c186 bl_186 br_186 wl_49 vdd gnd cell_6t
Xbit_r50_c186 bl_186 br_186 wl_50 vdd gnd cell_6t
Xbit_r51_c186 bl_186 br_186 wl_51 vdd gnd cell_6t
Xbit_r52_c186 bl_186 br_186 wl_52 vdd gnd cell_6t
Xbit_r53_c186 bl_186 br_186 wl_53 vdd gnd cell_6t
Xbit_r54_c186 bl_186 br_186 wl_54 vdd gnd cell_6t
Xbit_r55_c186 bl_186 br_186 wl_55 vdd gnd cell_6t
Xbit_r56_c186 bl_186 br_186 wl_56 vdd gnd cell_6t
Xbit_r57_c186 bl_186 br_186 wl_57 vdd gnd cell_6t
Xbit_r58_c186 bl_186 br_186 wl_58 vdd gnd cell_6t
Xbit_r59_c186 bl_186 br_186 wl_59 vdd gnd cell_6t
Xbit_r60_c186 bl_186 br_186 wl_60 vdd gnd cell_6t
Xbit_r61_c186 bl_186 br_186 wl_61 vdd gnd cell_6t
Xbit_r62_c186 bl_186 br_186 wl_62 vdd gnd cell_6t
Xbit_r63_c186 bl_186 br_186 wl_63 vdd gnd cell_6t
Xbit_r64_c186 bl_186 br_186 wl_64 vdd gnd cell_6t
Xbit_r65_c186 bl_186 br_186 wl_65 vdd gnd cell_6t
Xbit_r66_c186 bl_186 br_186 wl_66 vdd gnd cell_6t
Xbit_r67_c186 bl_186 br_186 wl_67 vdd gnd cell_6t
Xbit_r68_c186 bl_186 br_186 wl_68 vdd gnd cell_6t
Xbit_r69_c186 bl_186 br_186 wl_69 vdd gnd cell_6t
Xbit_r70_c186 bl_186 br_186 wl_70 vdd gnd cell_6t
Xbit_r71_c186 bl_186 br_186 wl_71 vdd gnd cell_6t
Xbit_r72_c186 bl_186 br_186 wl_72 vdd gnd cell_6t
Xbit_r73_c186 bl_186 br_186 wl_73 vdd gnd cell_6t
Xbit_r74_c186 bl_186 br_186 wl_74 vdd gnd cell_6t
Xbit_r75_c186 bl_186 br_186 wl_75 vdd gnd cell_6t
Xbit_r76_c186 bl_186 br_186 wl_76 vdd gnd cell_6t
Xbit_r77_c186 bl_186 br_186 wl_77 vdd gnd cell_6t
Xbit_r78_c186 bl_186 br_186 wl_78 vdd gnd cell_6t
Xbit_r79_c186 bl_186 br_186 wl_79 vdd gnd cell_6t
Xbit_r80_c186 bl_186 br_186 wl_80 vdd gnd cell_6t
Xbit_r81_c186 bl_186 br_186 wl_81 vdd gnd cell_6t
Xbit_r82_c186 bl_186 br_186 wl_82 vdd gnd cell_6t
Xbit_r83_c186 bl_186 br_186 wl_83 vdd gnd cell_6t
Xbit_r84_c186 bl_186 br_186 wl_84 vdd gnd cell_6t
Xbit_r85_c186 bl_186 br_186 wl_85 vdd gnd cell_6t
Xbit_r86_c186 bl_186 br_186 wl_86 vdd gnd cell_6t
Xbit_r87_c186 bl_186 br_186 wl_87 vdd gnd cell_6t
Xbit_r88_c186 bl_186 br_186 wl_88 vdd gnd cell_6t
Xbit_r89_c186 bl_186 br_186 wl_89 vdd gnd cell_6t
Xbit_r90_c186 bl_186 br_186 wl_90 vdd gnd cell_6t
Xbit_r91_c186 bl_186 br_186 wl_91 vdd gnd cell_6t
Xbit_r92_c186 bl_186 br_186 wl_92 vdd gnd cell_6t
Xbit_r93_c186 bl_186 br_186 wl_93 vdd gnd cell_6t
Xbit_r94_c186 bl_186 br_186 wl_94 vdd gnd cell_6t
Xbit_r95_c186 bl_186 br_186 wl_95 vdd gnd cell_6t
Xbit_r96_c186 bl_186 br_186 wl_96 vdd gnd cell_6t
Xbit_r97_c186 bl_186 br_186 wl_97 vdd gnd cell_6t
Xbit_r98_c186 bl_186 br_186 wl_98 vdd gnd cell_6t
Xbit_r99_c186 bl_186 br_186 wl_99 vdd gnd cell_6t
Xbit_r100_c186 bl_186 br_186 wl_100 vdd gnd cell_6t
Xbit_r101_c186 bl_186 br_186 wl_101 vdd gnd cell_6t
Xbit_r102_c186 bl_186 br_186 wl_102 vdd gnd cell_6t
Xbit_r103_c186 bl_186 br_186 wl_103 vdd gnd cell_6t
Xbit_r104_c186 bl_186 br_186 wl_104 vdd gnd cell_6t
Xbit_r105_c186 bl_186 br_186 wl_105 vdd gnd cell_6t
Xbit_r106_c186 bl_186 br_186 wl_106 vdd gnd cell_6t
Xbit_r107_c186 bl_186 br_186 wl_107 vdd gnd cell_6t
Xbit_r108_c186 bl_186 br_186 wl_108 vdd gnd cell_6t
Xbit_r109_c186 bl_186 br_186 wl_109 vdd gnd cell_6t
Xbit_r110_c186 bl_186 br_186 wl_110 vdd gnd cell_6t
Xbit_r111_c186 bl_186 br_186 wl_111 vdd gnd cell_6t
Xbit_r112_c186 bl_186 br_186 wl_112 vdd gnd cell_6t
Xbit_r113_c186 bl_186 br_186 wl_113 vdd gnd cell_6t
Xbit_r114_c186 bl_186 br_186 wl_114 vdd gnd cell_6t
Xbit_r115_c186 bl_186 br_186 wl_115 vdd gnd cell_6t
Xbit_r116_c186 bl_186 br_186 wl_116 vdd gnd cell_6t
Xbit_r117_c186 bl_186 br_186 wl_117 vdd gnd cell_6t
Xbit_r118_c186 bl_186 br_186 wl_118 vdd gnd cell_6t
Xbit_r119_c186 bl_186 br_186 wl_119 vdd gnd cell_6t
Xbit_r120_c186 bl_186 br_186 wl_120 vdd gnd cell_6t
Xbit_r121_c186 bl_186 br_186 wl_121 vdd gnd cell_6t
Xbit_r122_c186 bl_186 br_186 wl_122 vdd gnd cell_6t
Xbit_r123_c186 bl_186 br_186 wl_123 vdd gnd cell_6t
Xbit_r124_c186 bl_186 br_186 wl_124 vdd gnd cell_6t
Xbit_r125_c186 bl_186 br_186 wl_125 vdd gnd cell_6t
Xbit_r126_c186 bl_186 br_186 wl_126 vdd gnd cell_6t
Xbit_r127_c186 bl_186 br_186 wl_127 vdd gnd cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd cell_6t
Xbit_r1_c187 bl_187 br_187 wl_1 vdd gnd cell_6t
Xbit_r2_c187 bl_187 br_187 wl_2 vdd gnd cell_6t
Xbit_r3_c187 bl_187 br_187 wl_3 vdd gnd cell_6t
Xbit_r4_c187 bl_187 br_187 wl_4 vdd gnd cell_6t
Xbit_r5_c187 bl_187 br_187 wl_5 vdd gnd cell_6t
Xbit_r6_c187 bl_187 br_187 wl_6 vdd gnd cell_6t
Xbit_r7_c187 bl_187 br_187 wl_7 vdd gnd cell_6t
Xbit_r8_c187 bl_187 br_187 wl_8 vdd gnd cell_6t
Xbit_r9_c187 bl_187 br_187 wl_9 vdd gnd cell_6t
Xbit_r10_c187 bl_187 br_187 wl_10 vdd gnd cell_6t
Xbit_r11_c187 bl_187 br_187 wl_11 vdd gnd cell_6t
Xbit_r12_c187 bl_187 br_187 wl_12 vdd gnd cell_6t
Xbit_r13_c187 bl_187 br_187 wl_13 vdd gnd cell_6t
Xbit_r14_c187 bl_187 br_187 wl_14 vdd gnd cell_6t
Xbit_r15_c187 bl_187 br_187 wl_15 vdd gnd cell_6t
Xbit_r16_c187 bl_187 br_187 wl_16 vdd gnd cell_6t
Xbit_r17_c187 bl_187 br_187 wl_17 vdd gnd cell_6t
Xbit_r18_c187 bl_187 br_187 wl_18 vdd gnd cell_6t
Xbit_r19_c187 bl_187 br_187 wl_19 vdd gnd cell_6t
Xbit_r20_c187 bl_187 br_187 wl_20 vdd gnd cell_6t
Xbit_r21_c187 bl_187 br_187 wl_21 vdd gnd cell_6t
Xbit_r22_c187 bl_187 br_187 wl_22 vdd gnd cell_6t
Xbit_r23_c187 bl_187 br_187 wl_23 vdd gnd cell_6t
Xbit_r24_c187 bl_187 br_187 wl_24 vdd gnd cell_6t
Xbit_r25_c187 bl_187 br_187 wl_25 vdd gnd cell_6t
Xbit_r26_c187 bl_187 br_187 wl_26 vdd gnd cell_6t
Xbit_r27_c187 bl_187 br_187 wl_27 vdd gnd cell_6t
Xbit_r28_c187 bl_187 br_187 wl_28 vdd gnd cell_6t
Xbit_r29_c187 bl_187 br_187 wl_29 vdd gnd cell_6t
Xbit_r30_c187 bl_187 br_187 wl_30 vdd gnd cell_6t
Xbit_r31_c187 bl_187 br_187 wl_31 vdd gnd cell_6t
Xbit_r32_c187 bl_187 br_187 wl_32 vdd gnd cell_6t
Xbit_r33_c187 bl_187 br_187 wl_33 vdd gnd cell_6t
Xbit_r34_c187 bl_187 br_187 wl_34 vdd gnd cell_6t
Xbit_r35_c187 bl_187 br_187 wl_35 vdd gnd cell_6t
Xbit_r36_c187 bl_187 br_187 wl_36 vdd gnd cell_6t
Xbit_r37_c187 bl_187 br_187 wl_37 vdd gnd cell_6t
Xbit_r38_c187 bl_187 br_187 wl_38 vdd gnd cell_6t
Xbit_r39_c187 bl_187 br_187 wl_39 vdd gnd cell_6t
Xbit_r40_c187 bl_187 br_187 wl_40 vdd gnd cell_6t
Xbit_r41_c187 bl_187 br_187 wl_41 vdd gnd cell_6t
Xbit_r42_c187 bl_187 br_187 wl_42 vdd gnd cell_6t
Xbit_r43_c187 bl_187 br_187 wl_43 vdd gnd cell_6t
Xbit_r44_c187 bl_187 br_187 wl_44 vdd gnd cell_6t
Xbit_r45_c187 bl_187 br_187 wl_45 vdd gnd cell_6t
Xbit_r46_c187 bl_187 br_187 wl_46 vdd gnd cell_6t
Xbit_r47_c187 bl_187 br_187 wl_47 vdd gnd cell_6t
Xbit_r48_c187 bl_187 br_187 wl_48 vdd gnd cell_6t
Xbit_r49_c187 bl_187 br_187 wl_49 vdd gnd cell_6t
Xbit_r50_c187 bl_187 br_187 wl_50 vdd gnd cell_6t
Xbit_r51_c187 bl_187 br_187 wl_51 vdd gnd cell_6t
Xbit_r52_c187 bl_187 br_187 wl_52 vdd gnd cell_6t
Xbit_r53_c187 bl_187 br_187 wl_53 vdd gnd cell_6t
Xbit_r54_c187 bl_187 br_187 wl_54 vdd gnd cell_6t
Xbit_r55_c187 bl_187 br_187 wl_55 vdd gnd cell_6t
Xbit_r56_c187 bl_187 br_187 wl_56 vdd gnd cell_6t
Xbit_r57_c187 bl_187 br_187 wl_57 vdd gnd cell_6t
Xbit_r58_c187 bl_187 br_187 wl_58 vdd gnd cell_6t
Xbit_r59_c187 bl_187 br_187 wl_59 vdd gnd cell_6t
Xbit_r60_c187 bl_187 br_187 wl_60 vdd gnd cell_6t
Xbit_r61_c187 bl_187 br_187 wl_61 vdd gnd cell_6t
Xbit_r62_c187 bl_187 br_187 wl_62 vdd gnd cell_6t
Xbit_r63_c187 bl_187 br_187 wl_63 vdd gnd cell_6t
Xbit_r64_c187 bl_187 br_187 wl_64 vdd gnd cell_6t
Xbit_r65_c187 bl_187 br_187 wl_65 vdd gnd cell_6t
Xbit_r66_c187 bl_187 br_187 wl_66 vdd gnd cell_6t
Xbit_r67_c187 bl_187 br_187 wl_67 vdd gnd cell_6t
Xbit_r68_c187 bl_187 br_187 wl_68 vdd gnd cell_6t
Xbit_r69_c187 bl_187 br_187 wl_69 vdd gnd cell_6t
Xbit_r70_c187 bl_187 br_187 wl_70 vdd gnd cell_6t
Xbit_r71_c187 bl_187 br_187 wl_71 vdd gnd cell_6t
Xbit_r72_c187 bl_187 br_187 wl_72 vdd gnd cell_6t
Xbit_r73_c187 bl_187 br_187 wl_73 vdd gnd cell_6t
Xbit_r74_c187 bl_187 br_187 wl_74 vdd gnd cell_6t
Xbit_r75_c187 bl_187 br_187 wl_75 vdd gnd cell_6t
Xbit_r76_c187 bl_187 br_187 wl_76 vdd gnd cell_6t
Xbit_r77_c187 bl_187 br_187 wl_77 vdd gnd cell_6t
Xbit_r78_c187 bl_187 br_187 wl_78 vdd gnd cell_6t
Xbit_r79_c187 bl_187 br_187 wl_79 vdd gnd cell_6t
Xbit_r80_c187 bl_187 br_187 wl_80 vdd gnd cell_6t
Xbit_r81_c187 bl_187 br_187 wl_81 vdd gnd cell_6t
Xbit_r82_c187 bl_187 br_187 wl_82 vdd gnd cell_6t
Xbit_r83_c187 bl_187 br_187 wl_83 vdd gnd cell_6t
Xbit_r84_c187 bl_187 br_187 wl_84 vdd gnd cell_6t
Xbit_r85_c187 bl_187 br_187 wl_85 vdd gnd cell_6t
Xbit_r86_c187 bl_187 br_187 wl_86 vdd gnd cell_6t
Xbit_r87_c187 bl_187 br_187 wl_87 vdd gnd cell_6t
Xbit_r88_c187 bl_187 br_187 wl_88 vdd gnd cell_6t
Xbit_r89_c187 bl_187 br_187 wl_89 vdd gnd cell_6t
Xbit_r90_c187 bl_187 br_187 wl_90 vdd gnd cell_6t
Xbit_r91_c187 bl_187 br_187 wl_91 vdd gnd cell_6t
Xbit_r92_c187 bl_187 br_187 wl_92 vdd gnd cell_6t
Xbit_r93_c187 bl_187 br_187 wl_93 vdd gnd cell_6t
Xbit_r94_c187 bl_187 br_187 wl_94 vdd gnd cell_6t
Xbit_r95_c187 bl_187 br_187 wl_95 vdd gnd cell_6t
Xbit_r96_c187 bl_187 br_187 wl_96 vdd gnd cell_6t
Xbit_r97_c187 bl_187 br_187 wl_97 vdd gnd cell_6t
Xbit_r98_c187 bl_187 br_187 wl_98 vdd gnd cell_6t
Xbit_r99_c187 bl_187 br_187 wl_99 vdd gnd cell_6t
Xbit_r100_c187 bl_187 br_187 wl_100 vdd gnd cell_6t
Xbit_r101_c187 bl_187 br_187 wl_101 vdd gnd cell_6t
Xbit_r102_c187 bl_187 br_187 wl_102 vdd gnd cell_6t
Xbit_r103_c187 bl_187 br_187 wl_103 vdd gnd cell_6t
Xbit_r104_c187 bl_187 br_187 wl_104 vdd gnd cell_6t
Xbit_r105_c187 bl_187 br_187 wl_105 vdd gnd cell_6t
Xbit_r106_c187 bl_187 br_187 wl_106 vdd gnd cell_6t
Xbit_r107_c187 bl_187 br_187 wl_107 vdd gnd cell_6t
Xbit_r108_c187 bl_187 br_187 wl_108 vdd gnd cell_6t
Xbit_r109_c187 bl_187 br_187 wl_109 vdd gnd cell_6t
Xbit_r110_c187 bl_187 br_187 wl_110 vdd gnd cell_6t
Xbit_r111_c187 bl_187 br_187 wl_111 vdd gnd cell_6t
Xbit_r112_c187 bl_187 br_187 wl_112 vdd gnd cell_6t
Xbit_r113_c187 bl_187 br_187 wl_113 vdd gnd cell_6t
Xbit_r114_c187 bl_187 br_187 wl_114 vdd gnd cell_6t
Xbit_r115_c187 bl_187 br_187 wl_115 vdd gnd cell_6t
Xbit_r116_c187 bl_187 br_187 wl_116 vdd gnd cell_6t
Xbit_r117_c187 bl_187 br_187 wl_117 vdd gnd cell_6t
Xbit_r118_c187 bl_187 br_187 wl_118 vdd gnd cell_6t
Xbit_r119_c187 bl_187 br_187 wl_119 vdd gnd cell_6t
Xbit_r120_c187 bl_187 br_187 wl_120 vdd gnd cell_6t
Xbit_r121_c187 bl_187 br_187 wl_121 vdd gnd cell_6t
Xbit_r122_c187 bl_187 br_187 wl_122 vdd gnd cell_6t
Xbit_r123_c187 bl_187 br_187 wl_123 vdd gnd cell_6t
Xbit_r124_c187 bl_187 br_187 wl_124 vdd gnd cell_6t
Xbit_r125_c187 bl_187 br_187 wl_125 vdd gnd cell_6t
Xbit_r126_c187 bl_187 br_187 wl_126 vdd gnd cell_6t
Xbit_r127_c187 bl_187 br_187 wl_127 vdd gnd cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd cell_6t
Xbit_r1_c188 bl_188 br_188 wl_1 vdd gnd cell_6t
Xbit_r2_c188 bl_188 br_188 wl_2 vdd gnd cell_6t
Xbit_r3_c188 bl_188 br_188 wl_3 vdd gnd cell_6t
Xbit_r4_c188 bl_188 br_188 wl_4 vdd gnd cell_6t
Xbit_r5_c188 bl_188 br_188 wl_5 vdd gnd cell_6t
Xbit_r6_c188 bl_188 br_188 wl_6 vdd gnd cell_6t
Xbit_r7_c188 bl_188 br_188 wl_7 vdd gnd cell_6t
Xbit_r8_c188 bl_188 br_188 wl_8 vdd gnd cell_6t
Xbit_r9_c188 bl_188 br_188 wl_9 vdd gnd cell_6t
Xbit_r10_c188 bl_188 br_188 wl_10 vdd gnd cell_6t
Xbit_r11_c188 bl_188 br_188 wl_11 vdd gnd cell_6t
Xbit_r12_c188 bl_188 br_188 wl_12 vdd gnd cell_6t
Xbit_r13_c188 bl_188 br_188 wl_13 vdd gnd cell_6t
Xbit_r14_c188 bl_188 br_188 wl_14 vdd gnd cell_6t
Xbit_r15_c188 bl_188 br_188 wl_15 vdd gnd cell_6t
Xbit_r16_c188 bl_188 br_188 wl_16 vdd gnd cell_6t
Xbit_r17_c188 bl_188 br_188 wl_17 vdd gnd cell_6t
Xbit_r18_c188 bl_188 br_188 wl_18 vdd gnd cell_6t
Xbit_r19_c188 bl_188 br_188 wl_19 vdd gnd cell_6t
Xbit_r20_c188 bl_188 br_188 wl_20 vdd gnd cell_6t
Xbit_r21_c188 bl_188 br_188 wl_21 vdd gnd cell_6t
Xbit_r22_c188 bl_188 br_188 wl_22 vdd gnd cell_6t
Xbit_r23_c188 bl_188 br_188 wl_23 vdd gnd cell_6t
Xbit_r24_c188 bl_188 br_188 wl_24 vdd gnd cell_6t
Xbit_r25_c188 bl_188 br_188 wl_25 vdd gnd cell_6t
Xbit_r26_c188 bl_188 br_188 wl_26 vdd gnd cell_6t
Xbit_r27_c188 bl_188 br_188 wl_27 vdd gnd cell_6t
Xbit_r28_c188 bl_188 br_188 wl_28 vdd gnd cell_6t
Xbit_r29_c188 bl_188 br_188 wl_29 vdd gnd cell_6t
Xbit_r30_c188 bl_188 br_188 wl_30 vdd gnd cell_6t
Xbit_r31_c188 bl_188 br_188 wl_31 vdd gnd cell_6t
Xbit_r32_c188 bl_188 br_188 wl_32 vdd gnd cell_6t
Xbit_r33_c188 bl_188 br_188 wl_33 vdd gnd cell_6t
Xbit_r34_c188 bl_188 br_188 wl_34 vdd gnd cell_6t
Xbit_r35_c188 bl_188 br_188 wl_35 vdd gnd cell_6t
Xbit_r36_c188 bl_188 br_188 wl_36 vdd gnd cell_6t
Xbit_r37_c188 bl_188 br_188 wl_37 vdd gnd cell_6t
Xbit_r38_c188 bl_188 br_188 wl_38 vdd gnd cell_6t
Xbit_r39_c188 bl_188 br_188 wl_39 vdd gnd cell_6t
Xbit_r40_c188 bl_188 br_188 wl_40 vdd gnd cell_6t
Xbit_r41_c188 bl_188 br_188 wl_41 vdd gnd cell_6t
Xbit_r42_c188 bl_188 br_188 wl_42 vdd gnd cell_6t
Xbit_r43_c188 bl_188 br_188 wl_43 vdd gnd cell_6t
Xbit_r44_c188 bl_188 br_188 wl_44 vdd gnd cell_6t
Xbit_r45_c188 bl_188 br_188 wl_45 vdd gnd cell_6t
Xbit_r46_c188 bl_188 br_188 wl_46 vdd gnd cell_6t
Xbit_r47_c188 bl_188 br_188 wl_47 vdd gnd cell_6t
Xbit_r48_c188 bl_188 br_188 wl_48 vdd gnd cell_6t
Xbit_r49_c188 bl_188 br_188 wl_49 vdd gnd cell_6t
Xbit_r50_c188 bl_188 br_188 wl_50 vdd gnd cell_6t
Xbit_r51_c188 bl_188 br_188 wl_51 vdd gnd cell_6t
Xbit_r52_c188 bl_188 br_188 wl_52 vdd gnd cell_6t
Xbit_r53_c188 bl_188 br_188 wl_53 vdd gnd cell_6t
Xbit_r54_c188 bl_188 br_188 wl_54 vdd gnd cell_6t
Xbit_r55_c188 bl_188 br_188 wl_55 vdd gnd cell_6t
Xbit_r56_c188 bl_188 br_188 wl_56 vdd gnd cell_6t
Xbit_r57_c188 bl_188 br_188 wl_57 vdd gnd cell_6t
Xbit_r58_c188 bl_188 br_188 wl_58 vdd gnd cell_6t
Xbit_r59_c188 bl_188 br_188 wl_59 vdd gnd cell_6t
Xbit_r60_c188 bl_188 br_188 wl_60 vdd gnd cell_6t
Xbit_r61_c188 bl_188 br_188 wl_61 vdd gnd cell_6t
Xbit_r62_c188 bl_188 br_188 wl_62 vdd gnd cell_6t
Xbit_r63_c188 bl_188 br_188 wl_63 vdd gnd cell_6t
Xbit_r64_c188 bl_188 br_188 wl_64 vdd gnd cell_6t
Xbit_r65_c188 bl_188 br_188 wl_65 vdd gnd cell_6t
Xbit_r66_c188 bl_188 br_188 wl_66 vdd gnd cell_6t
Xbit_r67_c188 bl_188 br_188 wl_67 vdd gnd cell_6t
Xbit_r68_c188 bl_188 br_188 wl_68 vdd gnd cell_6t
Xbit_r69_c188 bl_188 br_188 wl_69 vdd gnd cell_6t
Xbit_r70_c188 bl_188 br_188 wl_70 vdd gnd cell_6t
Xbit_r71_c188 bl_188 br_188 wl_71 vdd gnd cell_6t
Xbit_r72_c188 bl_188 br_188 wl_72 vdd gnd cell_6t
Xbit_r73_c188 bl_188 br_188 wl_73 vdd gnd cell_6t
Xbit_r74_c188 bl_188 br_188 wl_74 vdd gnd cell_6t
Xbit_r75_c188 bl_188 br_188 wl_75 vdd gnd cell_6t
Xbit_r76_c188 bl_188 br_188 wl_76 vdd gnd cell_6t
Xbit_r77_c188 bl_188 br_188 wl_77 vdd gnd cell_6t
Xbit_r78_c188 bl_188 br_188 wl_78 vdd gnd cell_6t
Xbit_r79_c188 bl_188 br_188 wl_79 vdd gnd cell_6t
Xbit_r80_c188 bl_188 br_188 wl_80 vdd gnd cell_6t
Xbit_r81_c188 bl_188 br_188 wl_81 vdd gnd cell_6t
Xbit_r82_c188 bl_188 br_188 wl_82 vdd gnd cell_6t
Xbit_r83_c188 bl_188 br_188 wl_83 vdd gnd cell_6t
Xbit_r84_c188 bl_188 br_188 wl_84 vdd gnd cell_6t
Xbit_r85_c188 bl_188 br_188 wl_85 vdd gnd cell_6t
Xbit_r86_c188 bl_188 br_188 wl_86 vdd gnd cell_6t
Xbit_r87_c188 bl_188 br_188 wl_87 vdd gnd cell_6t
Xbit_r88_c188 bl_188 br_188 wl_88 vdd gnd cell_6t
Xbit_r89_c188 bl_188 br_188 wl_89 vdd gnd cell_6t
Xbit_r90_c188 bl_188 br_188 wl_90 vdd gnd cell_6t
Xbit_r91_c188 bl_188 br_188 wl_91 vdd gnd cell_6t
Xbit_r92_c188 bl_188 br_188 wl_92 vdd gnd cell_6t
Xbit_r93_c188 bl_188 br_188 wl_93 vdd gnd cell_6t
Xbit_r94_c188 bl_188 br_188 wl_94 vdd gnd cell_6t
Xbit_r95_c188 bl_188 br_188 wl_95 vdd gnd cell_6t
Xbit_r96_c188 bl_188 br_188 wl_96 vdd gnd cell_6t
Xbit_r97_c188 bl_188 br_188 wl_97 vdd gnd cell_6t
Xbit_r98_c188 bl_188 br_188 wl_98 vdd gnd cell_6t
Xbit_r99_c188 bl_188 br_188 wl_99 vdd gnd cell_6t
Xbit_r100_c188 bl_188 br_188 wl_100 vdd gnd cell_6t
Xbit_r101_c188 bl_188 br_188 wl_101 vdd gnd cell_6t
Xbit_r102_c188 bl_188 br_188 wl_102 vdd gnd cell_6t
Xbit_r103_c188 bl_188 br_188 wl_103 vdd gnd cell_6t
Xbit_r104_c188 bl_188 br_188 wl_104 vdd gnd cell_6t
Xbit_r105_c188 bl_188 br_188 wl_105 vdd gnd cell_6t
Xbit_r106_c188 bl_188 br_188 wl_106 vdd gnd cell_6t
Xbit_r107_c188 bl_188 br_188 wl_107 vdd gnd cell_6t
Xbit_r108_c188 bl_188 br_188 wl_108 vdd gnd cell_6t
Xbit_r109_c188 bl_188 br_188 wl_109 vdd gnd cell_6t
Xbit_r110_c188 bl_188 br_188 wl_110 vdd gnd cell_6t
Xbit_r111_c188 bl_188 br_188 wl_111 vdd gnd cell_6t
Xbit_r112_c188 bl_188 br_188 wl_112 vdd gnd cell_6t
Xbit_r113_c188 bl_188 br_188 wl_113 vdd gnd cell_6t
Xbit_r114_c188 bl_188 br_188 wl_114 vdd gnd cell_6t
Xbit_r115_c188 bl_188 br_188 wl_115 vdd gnd cell_6t
Xbit_r116_c188 bl_188 br_188 wl_116 vdd gnd cell_6t
Xbit_r117_c188 bl_188 br_188 wl_117 vdd gnd cell_6t
Xbit_r118_c188 bl_188 br_188 wl_118 vdd gnd cell_6t
Xbit_r119_c188 bl_188 br_188 wl_119 vdd gnd cell_6t
Xbit_r120_c188 bl_188 br_188 wl_120 vdd gnd cell_6t
Xbit_r121_c188 bl_188 br_188 wl_121 vdd gnd cell_6t
Xbit_r122_c188 bl_188 br_188 wl_122 vdd gnd cell_6t
Xbit_r123_c188 bl_188 br_188 wl_123 vdd gnd cell_6t
Xbit_r124_c188 bl_188 br_188 wl_124 vdd gnd cell_6t
Xbit_r125_c188 bl_188 br_188 wl_125 vdd gnd cell_6t
Xbit_r126_c188 bl_188 br_188 wl_126 vdd gnd cell_6t
Xbit_r127_c188 bl_188 br_188 wl_127 vdd gnd cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd cell_6t
Xbit_r1_c189 bl_189 br_189 wl_1 vdd gnd cell_6t
Xbit_r2_c189 bl_189 br_189 wl_2 vdd gnd cell_6t
Xbit_r3_c189 bl_189 br_189 wl_3 vdd gnd cell_6t
Xbit_r4_c189 bl_189 br_189 wl_4 vdd gnd cell_6t
Xbit_r5_c189 bl_189 br_189 wl_5 vdd gnd cell_6t
Xbit_r6_c189 bl_189 br_189 wl_6 vdd gnd cell_6t
Xbit_r7_c189 bl_189 br_189 wl_7 vdd gnd cell_6t
Xbit_r8_c189 bl_189 br_189 wl_8 vdd gnd cell_6t
Xbit_r9_c189 bl_189 br_189 wl_9 vdd gnd cell_6t
Xbit_r10_c189 bl_189 br_189 wl_10 vdd gnd cell_6t
Xbit_r11_c189 bl_189 br_189 wl_11 vdd gnd cell_6t
Xbit_r12_c189 bl_189 br_189 wl_12 vdd gnd cell_6t
Xbit_r13_c189 bl_189 br_189 wl_13 vdd gnd cell_6t
Xbit_r14_c189 bl_189 br_189 wl_14 vdd gnd cell_6t
Xbit_r15_c189 bl_189 br_189 wl_15 vdd gnd cell_6t
Xbit_r16_c189 bl_189 br_189 wl_16 vdd gnd cell_6t
Xbit_r17_c189 bl_189 br_189 wl_17 vdd gnd cell_6t
Xbit_r18_c189 bl_189 br_189 wl_18 vdd gnd cell_6t
Xbit_r19_c189 bl_189 br_189 wl_19 vdd gnd cell_6t
Xbit_r20_c189 bl_189 br_189 wl_20 vdd gnd cell_6t
Xbit_r21_c189 bl_189 br_189 wl_21 vdd gnd cell_6t
Xbit_r22_c189 bl_189 br_189 wl_22 vdd gnd cell_6t
Xbit_r23_c189 bl_189 br_189 wl_23 vdd gnd cell_6t
Xbit_r24_c189 bl_189 br_189 wl_24 vdd gnd cell_6t
Xbit_r25_c189 bl_189 br_189 wl_25 vdd gnd cell_6t
Xbit_r26_c189 bl_189 br_189 wl_26 vdd gnd cell_6t
Xbit_r27_c189 bl_189 br_189 wl_27 vdd gnd cell_6t
Xbit_r28_c189 bl_189 br_189 wl_28 vdd gnd cell_6t
Xbit_r29_c189 bl_189 br_189 wl_29 vdd gnd cell_6t
Xbit_r30_c189 bl_189 br_189 wl_30 vdd gnd cell_6t
Xbit_r31_c189 bl_189 br_189 wl_31 vdd gnd cell_6t
Xbit_r32_c189 bl_189 br_189 wl_32 vdd gnd cell_6t
Xbit_r33_c189 bl_189 br_189 wl_33 vdd gnd cell_6t
Xbit_r34_c189 bl_189 br_189 wl_34 vdd gnd cell_6t
Xbit_r35_c189 bl_189 br_189 wl_35 vdd gnd cell_6t
Xbit_r36_c189 bl_189 br_189 wl_36 vdd gnd cell_6t
Xbit_r37_c189 bl_189 br_189 wl_37 vdd gnd cell_6t
Xbit_r38_c189 bl_189 br_189 wl_38 vdd gnd cell_6t
Xbit_r39_c189 bl_189 br_189 wl_39 vdd gnd cell_6t
Xbit_r40_c189 bl_189 br_189 wl_40 vdd gnd cell_6t
Xbit_r41_c189 bl_189 br_189 wl_41 vdd gnd cell_6t
Xbit_r42_c189 bl_189 br_189 wl_42 vdd gnd cell_6t
Xbit_r43_c189 bl_189 br_189 wl_43 vdd gnd cell_6t
Xbit_r44_c189 bl_189 br_189 wl_44 vdd gnd cell_6t
Xbit_r45_c189 bl_189 br_189 wl_45 vdd gnd cell_6t
Xbit_r46_c189 bl_189 br_189 wl_46 vdd gnd cell_6t
Xbit_r47_c189 bl_189 br_189 wl_47 vdd gnd cell_6t
Xbit_r48_c189 bl_189 br_189 wl_48 vdd gnd cell_6t
Xbit_r49_c189 bl_189 br_189 wl_49 vdd gnd cell_6t
Xbit_r50_c189 bl_189 br_189 wl_50 vdd gnd cell_6t
Xbit_r51_c189 bl_189 br_189 wl_51 vdd gnd cell_6t
Xbit_r52_c189 bl_189 br_189 wl_52 vdd gnd cell_6t
Xbit_r53_c189 bl_189 br_189 wl_53 vdd gnd cell_6t
Xbit_r54_c189 bl_189 br_189 wl_54 vdd gnd cell_6t
Xbit_r55_c189 bl_189 br_189 wl_55 vdd gnd cell_6t
Xbit_r56_c189 bl_189 br_189 wl_56 vdd gnd cell_6t
Xbit_r57_c189 bl_189 br_189 wl_57 vdd gnd cell_6t
Xbit_r58_c189 bl_189 br_189 wl_58 vdd gnd cell_6t
Xbit_r59_c189 bl_189 br_189 wl_59 vdd gnd cell_6t
Xbit_r60_c189 bl_189 br_189 wl_60 vdd gnd cell_6t
Xbit_r61_c189 bl_189 br_189 wl_61 vdd gnd cell_6t
Xbit_r62_c189 bl_189 br_189 wl_62 vdd gnd cell_6t
Xbit_r63_c189 bl_189 br_189 wl_63 vdd gnd cell_6t
Xbit_r64_c189 bl_189 br_189 wl_64 vdd gnd cell_6t
Xbit_r65_c189 bl_189 br_189 wl_65 vdd gnd cell_6t
Xbit_r66_c189 bl_189 br_189 wl_66 vdd gnd cell_6t
Xbit_r67_c189 bl_189 br_189 wl_67 vdd gnd cell_6t
Xbit_r68_c189 bl_189 br_189 wl_68 vdd gnd cell_6t
Xbit_r69_c189 bl_189 br_189 wl_69 vdd gnd cell_6t
Xbit_r70_c189 bl_189 br_189 wl_70 vdd gnd cell_6t
Xbit_r71_c189 bl_189 br_189 wl_71 vdd gnd cell_6t
Xbit_r72_c189 bl_189 br_189 wl_72 vdd gnd cell_6t
Xbit_r73_c189 bl_189 br_189 wl_73 vdd gnd cell_6t
Xbit_r74_c189 bl_189 br_189 wl_74 vdd gnd cell_6t
Xbit_r75_c189 bl_189 br_189 wl_75 vdd gnd cell_6t
Xbit_r76_c189 bl_189 br_189 wl_76 vdd gnd cell_6t
Xbit_r77_c189 bl_189 br_189 wl_77 vdd gnd cell_6t
Xbit_r78_c189 bl_189 br_189 wl_78 vdd gnd cell_6t
Xbit_r79_c189 bl_189 br_189 wl_79 vdd gnd cell_6t
Xbit_r80_c189 bl_189 br_189 wl_80 vdd gnd cell_6t
Xbit_r81_c189 bl_189 br_189 wl_81 vdd gnd cell_6t
Xbit_r82_c189 bl_189 br_189 wl_82 vdd gnd cell_6t
Xbit_r83_c189 bl_189 br_189 wl_83 vdd gnd cell_6t
Xbit_r84_c189 bl_189 br_189 wl_84 vdd gnd cell_6t
Xbit_r85_c189 bl_189 br_189 wl_85 vdd gnd cell_6t
Xbit_r86_c189 bl_189 br_189 wl_86 vdd gnd cell_6t
Xbit_r87_c189 bl_189 br_189 wl_87 vdd gnd cell_6t
Xbit_r88_c189 bl_189 br_189 wl_88 vdd gnd cell_6t
Xbit_r89_c189 bl_189 br_189 wl_89 vdd gnd cell_6t
Xbit_r90_c189 bl_189 br_189 wl_90 vdd gnd cell_6t
Xbit_r91_c189 bl_189 br_189 wl_91 vdd gnd cell_6t
Xbit_r92_c189 bl_189 br_189 wl_92 vdd gnd cell_6t
Xbit_r93_c189 bl_189 br_189 wl_93 vdd gnd cell_6t
Xbit_r94_c189 bl_189 br_189 wl_94 vdd gnd cell_6t
Xbit_r95_c189 bl_189 br_189 wl_95 vdd gnd cell_6t
Xbit_r96_c189 bl_189 br_189 wl_96 vdd gnd cell_6t
Xbit_r97_c189 bl_189 br_189 wl_97 vdd gnd cell_6t
Xbit_r98_c189 bl_189 br_189 wl_98 vdd gnd cell_6t
Xbit_r99_c189 bl_189 br_189 wl_99 vdd gnd cell_6t
Xbit_r100_c189 bl_189 br_189 wl_100 vdd gnd cell_6t
Xbit_r101_c189 bl_189 br_189 wl_101 vdd gnd cell_6t
Xbit_r102_c189 bl_189 br_189 wl_102 vdd gnd cell_6t
Xbit_r103_c189 bl_189 br_189 wl_103 vdd gnd cell_6t
Xbit_r104_c189 bl_189 br_189 wl_104 vdd gnd cell_6t
Xbit_r105_c189 bl_189 br_189 wl_105 vdd gnd cell_6t
Xbit_r106_c189 bl_189 br_189 wl_106 vdd gnd cell_6t
Xbit_r107_c189 bl_189 br_189 wl_107 vdd gnd cell_6t
Xbit_r108_c189 bl_189 br_189 wl_108 vdd gnd cell_6t
Xbit_r109_c189 bl_189 br_189 wl_109 vdd gnd cell_6t
Xbit_r110_c189 bl_189 br_189 wl_110 vdd gnd cell_6t
Xbit_r111_c189 bl_189 br_189 wl_111 vdd gnd cell_6t
Xbit_r112_c189 bl_189 br_189 wl_112 vdd gnd cell_6t
Xbit_r113_c189 bl_189 br_189 wl_113 vdd gnd cell_6t
Xbit_r114_c189 bl_189 br_189 wl_114 vdd gnd cell_6t
Xbit_r115_c189 bl_189 br_189 wl_115 vdd gnd cell_6t
Xbit_r116_c189 bl_189 br_189 wl_116 vdd gnd cell_6t
Xbit_r117_c189 bl_189 br_189 wl_117 vdd gnd cell_6t
Xbit_r118_c189 bl_189 br_189 wl_118 vdd gnd cell_6t
Xbit_r119_c189 bl_189 br_189 wl_119 vdd gnd cell_6t
Xbit_r120_c189 bl_189 br_189 wl_120 vdd gnd cell_6t
Xbit_r121_c189 bl_189 br_189 wl_121 vdd gnd cell_6t
Xbit_r122_c189 bl_189 br_189 wl_122 vdd gnd cell_6t
Xbit_r123_c189 bl_189 br_189 wl_123 vdd gnd cell_6t
Xbit_r124_c189 bl_189 br_189 wl_124 vdd gnd cell_6t
Xbit_r125_c189 bl_189 br_189 wl_125 vdd gnd cell_6t
Xbit_r126_c189 bl_189 br_189 wl_126 vdd gnd cell_6t
Xbit_r127_c189 bl_189 br_189 wl_127 vdd gnd cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd cell_6t
Xbit_r1_c190 bl_190 br_190 wl_1 vdd gnd cell_6t
Xbit_r2_c190 bl_190 br_190 wl_2 vdd gnd cell_6t
Xbit_r3_c190 bl_190 br_190 wl_3 vdd gnd cell_6t
Xbit_r4_c190 bl_190 br_190 wl_4 vdd gnd cell_6t
Xbit_r5_c190 bl_190 br_190 wl_5 vdd gnd cell_6t
Xbit_r6_c190 bl_190 br_190 wl_6 vdd gnd cell_6t
Xbit_r7_c190 bl_190 br_190 wl_7 vdd gnd cell_6t
Xbit_r8_c190 bl_190 br_190 wl_8 vdd gnd cell_6t
Xbit_r9_c190 bl_190 br_190 wl_9 vdd gnd cell_6t
Xbit_r10_c190 bl_190 br_190 wl_10 vdd gnd cell_6t
Xbit_r11_c190 bl_190 br_190 wl_11 vdd gnd cell_6t
Xbit_r12_c190 bl_190 br_190 wl_12 vdd gnd cell_6t
Xbit_r13_c190 bl_190 br_190 wl_13 vdd gnd cell_6t
Xbit_r14_c190 bl_190 br_190 wl_14 vdd gnd cell_6t
Xbit_r15_c190 bl_190 br_190 wl_15 vdd gnd cell_6t
Xbit_r16_c190 bl_190 br_190 wl_16 vdd gnd cell_6t
Xbit_r17_c190 bl_190 br_190 wl_17 vdd gnd cell_6t
Xbit_r18_c190 bl_190 br_190 wl_18 vdd gnd cell_6t
Xbit_r19_c190 bl_190 br_190 wl_19 vdd gnd cell_6t
Xbit_r20_c190 bl_190 br_190 wl_20 vdd gnd cell_6t
Xbit_r21_c190 bl_190 br_190 wl_21 vdd gnd cell_6t
Xbit_r22_c190 bl_190 br_190 wl_22 vdd gnd cell_6t
Xbit_r23_c190 bl_190 br_190 wl_23 vdd gnd cell_6t
Xbit_r24_c190 bl_190 br_190 wl_24 vdd gnd cell_6t
Xbit_r25_c190 bl_190 br_190 wl_25 vdd gnd cell_6t
Xbit_r26_c190 bl_190 br_190 wl_26 vdd gnd cell_6t
Xbit_r27_c190 bl_190 br_190 wl_27 vdd gnd cell_6t
Xbit_r28_c190 bl_190 br_190 wl_28 vdd gnd cell_6t
Xbit_r29_c190 bl_190 br_190 wl_29 vdd gnd cell_6t
Xbit_r30_c190 bl_190 br_190 wl_30 vdd gnd cell_6t
Xbit_r31_c190 bl_190 br_190 wl_31 vdd gnd cell_6t
Xbit_r32_c190 bl_190 br_190 wl_32 vdd gnd cell_6t
Xbit_r33_c190 bl_190 br_190 wl_33 vdd gnd cell_6t
Xbit_r34_c190 bl_190 br_190 wl_34 vdd gnd cell_6t
Xbit_r35_c190 bl_190 br_190 wl_35 vdd gnd cell_6t
Xbit_r36_c190 bl_190 br_190 wl_36 vdd gnd cell_6t
Xbit_r37_c190 bl_190 br_190 wl_37 vdd gnd cell_6t
Xbit_r38_c190 bl_190 br_190 wl_38 vdd gnd cell_6t
Xbit_r39_c190 bl_190 br_190 wl_39 vdd gnd cell_6t
Xbit_r40_c190 bl_190 br_190 wl_40 vdd gnd cell_6t
Xbit_r41_c190 bl_190 br_190 wl_41 vdd gnd cell_6t
Xbit_r42_c190 bl_190 br_190 wl_42 vdd gnd cell_6t
Xbit_r43_c190 bl_190 br_190 wl_43 vdd gnd cell_6t
Xbit_r44_c190 bl_190 br_190 wl_44 vdd gnd cell_6t
Xbit_r45_c190 bl_190 br_190 wl_45 vdd gnd cell_6t
Xbit_r46_c190 bl_190 br_190 wl_46 vdd gnd cell_6t
Xbit_r47_c190 bl_190 br_190 wl_47 vdd gnd cell_6t
Xbit_r48_c190 bl_190 br_190 wl_48 vdd gnd cell_6t
Xbit_r49_c190 bl_190 br_190 wl_49 vdd gnd cell_6t
Xbit_r50_c190 bl_190 br_190 wl_50 vdd gnd cell_6t
Xbit_r51_c190 bl_190 br_190 wl_51 vdd gnd cell_6t
Xbit_r52_c190 bl_190 br_190 wl_52 vdd gnd cell_6t
Xbit_r53_c190 bl_190 br_190 wl_53 vdd gnd cell_6t
Xbit_r54_c190 bl_190 br_190 wl_54 vdd gnd cell_6t
Xbit_r55_c190 bl_190 br_190 wl_55 vdd gnd cell_6t
Xbit_r56_c190 bl_190 br_190 wl_56 vdd gnd cell_6t
Xbit_r57_c190 bl_190 br_190 wl_57 vdd gnd cell_6t
Xbit_r58_c190 bl_190 br_190 wl_58 vdd gnd cell_6t
Xbit_r59_c190 bl_190 br_190 wl_59 vdd gnd cell_6t
Xbit_r60_c190 bl_190 br_190 wl_60 vdd gnd cell_6t
Xbit_r61_c190 bl_190 br_190 wl_61 vdd gnd cell_6t
Xbit_r62_c190 bl_190 br_190 wl_62 vdd gnd cell_6t
Xbit_r63_c190 bl_190 br_190 wl_63 vdd gnd cell_6t
Xbit_r64_c190 bl_190 br_190 wl_64 vdd gnd cell_6t
Xbit_r65_c190 bl_190 br_190 wl_65 vdd gnd cell_6t
Xbit_r66_c190 bl_190 br_190 wl_66 vdd gnd cell_6t
Xbit_r67_c190 bl_190 br_190 wl_67 vdd gnd cell_6t
Xbit_r68_c190 bl_190 br_190 wl_68 vdd gnd cell_6t
Xbit_r69_c190 bl_190 br_190 wl_69 vdd gnd cell_6t
Xbit_r70_c190 bl_190 br_190 wl_70 vdd gnd cell_6t
Xbit_r71_c190 bl_190 br_190 wl_71 vdd gnd cell_6t
Xbit_r72_c190 bl_190 br_190 wl_72 vdd gnd cell_6t
Xbit_r73_c190 bl_190 br_190 wl_73 vdd gnd cell_6t
Xbit_r74_c190 bl_190 br_190 wl_74 vdd gnd cell_6t
Xbit_r75_c190 bl_190 br_190 wl_75 vdd gnd cell_6t
Xbit_r76_c190 bl_190 br_190 wl_76 vdd gnd cell_6t
Xbit_r77_c190 bl_190 br_190 wl_77 vdd gnd cell_6t
Xbit_r78_c190 bl_190 br_190 wl_78 vdd gnd cell_6t
Xbit_r79_c190 bl_190 br_190 wl_79 vdd gnd cell_6t
Xbit_r80_c190 bl_190 br_190 wl_80 vdd gnd cell_6t
Xbit_r81_c190 bl_190 br_190 wl_81 vdd gnd cell_6t
Xbit_r82_c190 bl_190 br_190 wl_82 vdd gnd cell_6t
Xbit_r83_c190 bl_190 br_190 wl_83 vdd gnd cell_6t
Xbit_r84_c190 bl_190 br_190 wl_84 vdd gnd cell_6t
Xbit_r85_c190 bl_190 br_190 wl_85 vdd gnd cell_6t
Xbit_r86_c190 bl_190 br_190 wl_86 vdd gnd cell_6t
Xbit_r87_c190 bl_190 br_190 wl_87 vdd gnd cell_6t
Xbit_r88_c190 bl_190 br_190 wl_88 vdd gnd cell_6t
Xbit_r89_c190 bl_190 br_190 wl_89 vdd gnd cell_6t
Xbit_r90_c190 bl_190 br_190 wl_90 vdd gnd cell_6t
Xbit_r91_c190 bl_190 br_190 wl_91 vdd gnd cell_6t
Xbit_r92_c190 bl_190 br_190 wl_92 vdd gnd cell_6t
Xbit_r93_c190 bl_190 br_190 wl_93 vdd gnd cell_6t
Xbit_r94_c190 bl_190 br_190 wl_94 vdd gnd cell_6t
Xbit_r95_c190 bl_190 br_190 wl_95 vdd gnd cell_6t
Xbit_r96_c190 bl_190 br_190 wl_96 vdd gnd cell_6t
Xbit_r97_c190 bl_190 br_190 wl_97 vdd gnd cell_6t
Xbit_r98_c190 bl_190 br_190 wl_98 vdd gnd cell_6t
Xbit_r99_c190 bl_190 br_190 wl_99 vdd gnd cell_6t
Xbit_r100_c190 bl_190 br_190 wl_100 vdd gnd cell_6t
Xbit_r101_c190 bl_190 br_190 wl_101 vdd gnd cell_6t
Xbit_r102_c190 bl_190 br_190 wl_102 vdd gnd cell_6t
Xbit_r103_c190 bl_190 br_190 wl_103 vdd gnd cell_6t
Xbit_r104_c190 bl_190 br_190 wl_104 vdd gnd cell_6t
Xbit_r105_c190 bl_190 br_190 wl_105 vdd gnd cell_6t
Xbit_r106_c190 bl_190 br_190 wl_106 vdd gnd cell_6t
Xbit_r107_c190 bl_190 br_190 wl_107 vdd gnd cell_6t
Xbit_r108_c190 bl_190 br_190 wl_108 vdd gnd cell_6t
Xbit_r109_c190 bl_190 br_190 wl_109 vdd gnd cell_6t
Xbit_r110_c190 bl_190 br_190 wl_110 vdd gnd cell_6t
Xbit_r111_c190 bl_190 br_190 wl_111 vdd gnd cell_6t
Xbit_r112_c190 bl_190 br_190 wl_112 vdd gnd cell_6t
Xbit_r113_c190 bl_190 br_190 wl_113 vdd gnd cell_6t
Xbit_r114_c190 bl_190 br_190 wl_114 vdd gnd cell_6t
Xbit_r115_c190 bl_190 br_190 wl_115 vdd gnd cell_6t
Xbit_r116_c190 bl_190 br_190 wl_116 vdd gnd cell_6t
Xbit_r117_c190 bl_190 br_190 wl_117 vdd gnd cell_6t
Xbit_r118_c190 bl_190 br_190 wl_118 vdd gnd cell_6t
Xbit_r119_c190 bl_190 br_190 wl_119 vdd gnd cell_6t
Xbit_r120_c190 bl_190 br_190 wl_120 vdd gnd cell_6t
Xbit_r121_c190 bl_190 br_190 wl_121 vdd gnd cell_6t
Xbit_r122_c190 bl_190 br_190 wl_122 vdd gnd cell_6t
Xbit_r123_c190 bl_190 br_190 wl_123 vdd gnd cell_6t
Xbit_r124_c190 bl_190 br_190 wl_124 vdd gnd cell_6t
Xbit_r125_c190 bl_190 br_190 wl_125 vdd gnd cell_6t
Xbit_r126_c190 bl_190 br_190 wl_126 vdd gnd cell_6t
Xbit_r127_c190 bl_190 br_190 wl_127 vdd gnd cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd cell_6t
Xbit_r1_c191 bl_191 br_191 wl_1 vdd gnd cell_6t
Xbit_r2_c191 bl_191 br_191 wl_2 vdd gnd cell_6t
Xbit_r3_c191 bl_191 br_191 wl_3 vdd gnd cell_6t
Xbit_r4_c191 bl_191 br_191 wl_4 vdd gnd cell_6t
Xbit_r5_c191 bl_191 br_191 wl_5 vdd gnd cell_6t
Xbit_r6_c191 bl_191 br_191 wl_6 vdd gnd cell_6t
Xbit_r7_c191 bl_191 br_191 wl_7 vdd gnd cell_6t
Xbit_r8_c191 bl_191 br_191 wl_8 vdd gnd cell_6t
Xbit_r9_c191 bl_191 br_191 wl_9 vdd gnd cell_6t
Xbit_r10_c191 bl_191 br_191 wl_10 vdd gnd cell_6t
Xbit_r11_c191 bl_191 br_191 wl_11 vdd gnd cell_6t
Xbit_r12_c191 bl_191 br_191 wl_12 vdd gnd cell_6t
Xbit_r13_c191 bl_191 br_191 wl_13 vdd gnd cell_6t
Xbit_r14_c191 bl_191 br_191 wl_14 vdd gnd cell_6t
Xbit_r15_c191 bl_191 br_191 wl_15 vdd gnd cell_6t
Xbit_r16_c191 bl_191 br_191 wl_16 vdd gnd cell_6t
Xbit_r17_c191 bl_191 br_191 wl_17 vdd gnd cell_6t
Xbit_r18_c191 bl_191 br_191 wl_18 vdd gnd cell_6t
Xbit_r19_c191 bl_191 br_191 wl_19 vdd gnd cell_6t
Xbit_r20_c191 bl_191 br_191 wl_20 vdd gnd cell_6t
Xbit_r21_c191 bl_191 br_191 wl_21 vdd gnd cell_6t
Xbit_r22_c191 bl_191 br_191 wl_22 vdd gnd cell_6t
Xbit_r23_c191 bl_191 br_191 wl_23 vdd gnd cell_6t
Xbit_r24_c191 bl_191 br_191 wl_24 vdd gnd cell_6t
Xbit_r25_c191 bl_191 br_191 wl_25 vdd gnd cell_6t
Xbit_r26_c191 bl_191 br_191 wl_26 vdd gnd cell_6t
Xbit_r27_c191 bl_191 br_191 wl_27 vdd gnd cell_6t
Xbit_r28_c191 bl_191 br_191 wl_28 vdd gnd cell_6t
Xbit_r29_c191 bl_191 br_191 wl_29 vdd gnd cell_6t
Xbit_r30_c191 bl_191 br_191 wl_30 vdd gnd cell_6t
Xbit_r31_c191 bl_191 br_191 wl_31 vdd gnd cell_6t
Xbit_r32_c191 bl_191 br_191 wl_32 vdd gnd cell_6t
Xbit_r33_c191 bl_191 br_191 wl_33 vdd gnd cell_6t
Xbit_r34_c191 bl_191 br_191 wl_34 vdd gnd cell_6t
Xbit_r35_c191 bl_191 br_191 wl_35 vdd gnd cell_6t
Xbit_r36_c191 bl_191 br_191 wl_36 vdd gnd cell_6t
Xbit_r37_c191 bl_191 br_191 wl_37 vdd gnd cell_6t
Xbit_r38_c191 bl_191 br_191 wl_38 vdd gnd cell_6t
Xbit_r39_c191 bl_191 br_191 wl_39 vdd gnd cell_6t
Xbit_r40_c191 bl_191 br_191 wl_40 vdd gnd cell_6t
Xbit_r41_c191 bl_191 br_191 wl_41 vdd gnd cell_6t
Xbit_r42_c191 bl_191 br_191 wl_42 vdd gnd cell_6t
Xbit_r43_c191 bl_191 br_191 wl_43 vdd gnd cell_6t
Xbit_r44_c191 bl_191 br_191 wl_44 vdd gnd cell_6t
Xbit_r45_c191 bl_191 br_191 wl_45 vdd gnd cell_6t
Xbit_r46_c191 bl_191 br_191 wl_46 vdd gnd cell_6t
Xbit_r47_c191 bl_191 br_191 wl_47 vdd gnd cell_6t
Xbit_r48_c191 bl_191 br_191 wl_48 vdd gnd cell_6t
Xbit_r49_c191 bl_191 br_191 wl_49 vdd gnd cell_6t
Xbit_r50_c191 bl_191 br_191 wl_50 vdd gnd cell_6t
Xbit_r51_c191 bl_191 br_191 wl_51 vdd gnd cell_6t
Xbit_r52_c191 bl_191 br_191 wl_52 vdd gnd cell_6t
Xbit_r53_c191 bl_191 br_191 wl_53 vdd gnd cell_6t
Xbit_r54_c191 bl_191 br_191 wl_54 vdd gnd cell_6t
Xbit_r55_c191 bl_191 br_191 wl_55 vdd gnd cell_6t
Xbit_r56_c191 bl_191 br_191 wl_56 vdd gnd cell_6t
Xbit_r57_c191 bl_191 br_191 wl_57 vdd gnd cell_6t
Xbit_r58_c191 bl_191 br_191 wl_58 vdd gnd cell_6t
Xbit_r59_c191 bl_191 br_191 wl_59 vdd gnd cell_6t
Xbit_r60_c191 bl_191 br_191 wl_60 vdd gnd cell_6t
Xbit_r61_c191 bl_191 br_191 wl_61 vdd gnd cell_6t
Xbit_r62_c191 bl_191 br_191 wl_62 vdd gnd cell_6t
Xbit_r63_c191 bl_191 br_191 wl_63 vdd gnd cell_6t
Xbit_r64_c191 bl_191 br_191 wl_64 vdd gnd cell_6t
Xbit_r65_c191 bl_191 br_191 wl_65 vdd gnd cell_6t
Xbit_r66_c191 bl_191 br_191 wl_66 vdd gnd cell_6t
Xbit_r67_c191 bl_191 br_191 wl_67 vdd gnd cell_6t
Xbit_r68_c191 bl_191 br_191 wl_68 vdd gnd cell_6t
Xbit_r69_c191 bl_191 br_191 wl_69 vdd gnd cell_6t
Xbit_r70_c191 bl_191 br_191 wl_70 vdd gnd cell_6t
Xbit_r71_c191 bl_191 br_191 wl_71 vdd gnd cell_6t
Xbit_r72_c191 bl_191 br_191 wl_72 vdd gnd cell_6t
Xbit_r73_c191 bl_191 br_191 wl_73 vdd gnd cell_6t
Xbit_r74_c191 bl_191 br_191 wl_74 vdd gnd cell_6t
Xbit_r75_c191 bl_191 br_191 wl_75 vdd gnd cell_6t
Xbit_r76_c191 bl_191 br_191 wl_76 vdd gnd cell_6t
Xbit_r77_c191 bl_191 br_191 wl_77 vdd gnd cell_6t
Xbit_r78_c191 bl_191 br_191 wl_78 vdd gnd cell_6t
Xbit_r79_c191 bl_191 br_191 wl_79 vdd gnd cell_6t
Xbit_r80_c191 bl_191 br_191 wl_80 vdd gnd cell_6t
Xbit_r81_c191 bl_191 br_191 wl_81 vdd gnd cell_6t
Xbit_r82_c191 bl_191 br_191 wl_82 vdd gnd cell_6t
Xbit_r83_c191 bl_191 br_191 wl_83 vdd gnd cell_6t
Xbit_r84_c191 bl_191 br_191 wl_84 vdd gnd cell_6t
Xbit_r85_c191 bl_191 br_191 wl_85 vdd gnd cell_6t
Xbit_r86_c191 bl_191 br_191 wl_86 vdd gnd cell_6t
Xbit_r87_c191 bl_191 br_191 wl_87 vdd gnd cell_6t
Xbit_r88_c191 bl_191 br_191 wl_88 vdd gnd cell_6t
Xbit_r89_c191 bl_191 br_191 wl_89 vdd gnd cell_6t
Xbit_r90_c191 bl_191 br_191 wl_90 vdd gnd cell_6t
Xbit_r91_c191 bl_191 br_191 wl_91 vdd gnd cell_6t
Xbit_r92_c191 bl_191 br_191 wl_92 vdd gnd cell_6t
Xbit_r93_c191 bl_191 br_191 wl_93 vdd gnd cell_6t
Xbit_r94_c191 bl_191 br_191 wl_94 vdd gnd cell_6t
Xbit_r95_c191 bl_191 br_191 wl_95 vdd gnd cell_6t
Xbit_r96_c191 bl_191 br_191 wl_96 vdd gnd cell_6t
Xbit_r97_c191 bl_191 br_191 wl_97 vdd gnd cell_6t
Xbit_r98_c191 bl_191 br_191 wl_98 vdd gnd cell_6t
Xbit_r99_c191 bl_191 br_191 wl_99 vdd gnd cell_6t
Xbit_r100_c191 bl_191 br_191 wl_100 vdd gnd cell_6t
Xbit_r101_c191 bl_191 br_191 wl_101 vdd gnd cell_6t
Xbit_r102_c191 bl_191 br_191 wl_102 vdd gnd cell_6t
Xbit_r103_c191 bl_191 br_191 wl_103 vdd gnd cell_6t
Xbit_r104_c191 bl_191 br_191 wl_104 vdd gnd cell_6t
Xbit_r105_c191 bl_191 br_191 wl_105 vdd gnd cell_6t
Xbit_r106_c191 bl_191 br_191 wl_106 vdd gnd cell_6t
Xbit_r107_c191 bl_191 br_191 wl_107 vdd gnd cell_6t
Xbit_r108_c191 bl_191 br_191 wl_108 vdd gnd cell_6t
Xbit_r109_c191 bl_191 br_191 wl_109 vdd gnd cell_6t
Xbit_r110_c191 bl_191 br_191 wl_110 vdd gnd cell_6t
Xbit_r111_c191 bl_191 br_191 wl_111 vdd gnd cell_6t
Xbit_r112_c191 bl_191 br_191 wl_112 vdd gnd cell_6t
Xbit_r113_c191 bl_191 br_191 wl_113 vdd gnd cell_6t
Xbit_r114_c191 bl_191 br_191 wl_114 vdd gnd cell_6t
Xbit_r115_c191 bl_191 br_191 wl_115 vdd gnd cell_6t
Xbit_r116_c191 bl_191 br_191 wl_116 vdd gnd cell_6t
Xbit_r117_c191 bl_191 br_191 wl_117 vdd gnd cell_6t
Xbit_r118_c191 bl_191 br_191 wl_118 vdd gnd cell_6t
Xbit_r119_c191 bl_191 br_191 wl_119 vdd gnd cell_6t
Xbit_r120_c191 bl_191 br_191 wl_120 vdd gnd cell_6t
Xbit_r121_c191 bl_191 br_191 wl_121 vdd gnd cell_6t
Xbit_r122_c191 bl_191 br_191 wl_122 vdd gnd cell_6t
Xbit_r123_c191 bl_191 br_191 wl_123 vdd gnd cell_6t
Xbit_r124_c191 bl_191 br_191 wl_124 vdd gnd cell_6t
Xbit_r125_c191 bl_191 br_191 wl_125 vdd gnd cell_6t
Xbit_r126_c191 bl_191 br_191 wl_126 vdd gnd cell_6t
Xbit_r127_c191 bl_191 br_191 wl_127 vdd gnd cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd cell_6t
Xbit_r1_c192 bl_192 br_192 wl_1 vdd gnd cell_6t
Xbit_r2_c192 bl_192 br_192 wl_2 vdd gnd cell_6t
Xbit_r3_c192 bl_192 br_192 wl_3 vdd gnd cell_6t
Xbit_r4_c192 bl_192 br_192 wl_4 vdd gnd cell_6t
Xbit_r5_c192 bl_192 br_192 wl_5 vdd gnd cell_6t
Xbit_r6_c192 bl_192 br_192 wl_6 vdd gnd cell_6t
Xbit_r7_c192 bl_192 br_192 wl_7 vdd gnd cell_6t
Xbit_r8_c192 bl_192 br_192 wl_8 vdd gnd cell_6t
Xbit_r9_c192 bl_192 br_192 wl_9 vdd gnd cell_6t
Xbit_r10_c192 bl_192 br_192 wl_10 vdd gnd cell_6t
Xbit_r11_c192 bl_192 br_192 wl_11 vdd gnd cell_6t
Xbit_r12_c192 bl_192 br_192 wl_12 vdd gnd cell_6t
Xbit_r13_c192 bl_192 br_192 wl_13 vdd gnd cell_6t
Xbit_r14_c192 bl_192 br_192 wl_14 vdd gnd cell_6t
Xbit_r15_c192 bl_192 br_192 wl_15 vdd gnd cell_6t
Xbit_r16_c192 bl_192 br_192 wl_16 vdd gnd cell_6t
Xbit_r17_c192 bl_192 br_192 wl_17 vdd gnd cell_6t
Xbit_r18_c192 bl_192 br_192 wl_18 vdd gnd cell_6t
Xbit_r19_c192 bl_192 br_192 wl_19 vdd gnd cell_6t
Xbit_r20_c192 bl_192 br_192 wl_20 vdd gnd cell_6t
Xbit_r21_c192 bl_192 br_192 wl_21 vdd gnd cell_6t
Xbit_r22_c192 bl_192 br_192 wl_22 vdd gnd cell_6t
Xbit_r23_c192 bl_192 br_192 wl_23 vdd gnd cell_6t
Xbit_r24_c192 bl_192 br_192 wl_24 vdd gnd cell_6t
Xbit_r25_c192 bl_192 br_192 wl_25 vdd gnd cell_6t
Xbit_r26_c192 bl_192 br_192 wl_26 vdd gnd cell_6t
Xbit_r27_c192 bl_192 br_192 wl_27 vdd gnd cell_6t
Xbit_r28_c192 bl_192 br_192 wl_28 vdd gnd cell_6t
Xbit_r29_c192 bl_192 br_192 wl_29 vdd gnd cell_6t
Xbit_r30_c192 bl_192 br_192 wl_30 vdd gnd cell_6t
Xbit_r31_c192 bl_192 br_192 wl_31 vdd gnd cell_6t
Xbit_r32_c192 bl_192 br_192 wl_32 vdd gnd cell_6t
Xbit_r33_c192 bl_192 br_192 wl_33 vdd gnd cell_6t
Xbit_r34_c192 bl_192 br_192 wl_34 vdd gnd cell_6t
Xbit_r35_c192 bl_192 br_192 wl_35 vdd gnd cell_6t
Xbit_r36_c192 bl_192 br_192 wl_36 vdd gnd cell_6t
Xbit_r37_c192 bl_192 br_192 wl_37 vdd gnd cell_6t
Xbit_r38_c192 bl_192 br_192 wl_38 vdd gnd cell_6t
Xbit_r39_c192 bl_192 br_192 wl_39 vdd gnd cell_6t
Xbit_r40_c192 bl_192 br_192 wl_40 vdd gnd cell_6t
Xbit_r41_c192 bl_192 br_192 wl_41 vdd gnd cell_6t
Xbit_r42_c192 bl_192 br_192 wl_42 vdd gnd cell_6t
Xbit_r43_c192 bl_192 br_192 wl_43 vdd gnd cell_6t
Xbit_r44_c192 bl_192 br_192 wl_44 vdd gnd cell_6t
Xbit_r45_c192 bl_192 br_192 wl_45 vdd gnd cell_6t
Xbit_r46_c192 bl_192 br_192 wl_46 vdd gnd cell_6t
Xbit_r47_c192 bl_192 br_192 wl_47 vdd gnd cell_6t
Xbit_r48_c192 bl_192 br_192 wl_48 vdd gnd cell_6t
Xbit_r49_c192 bl_192 br_192 wl_49 vdd gnd cell_6t
Xbit_r50_c192 bl_192 br_192 wl_50 vdd gnd cell_6t
Xbit_r51_c192 bl_192 br_192 wl_51 vdd gnd cell_6t
Xbit_r52_c192 bl_192 br_192 wl_52 vdd gnd cell_6t
Xbit_r53_c192 bl_192 br_192 wl_53 vdd gnd cell_6t
Xbit_r54_c192 bl_192 br_192 wl_54 vdd gnd cell_6t
Xbit_r55_c192 bl_192 br_192 wl_55 vdd gnd cell_6t
Xbit_r56_c192 bl_192 br_192 wl_56 vdd gnd cell_6t
Xbit_r57_c192 bl_192 br_192 wl_57 vdd gnd cell_6t
Xbit_r58_c192 bl_192 br_192 wl_58 vdd gnd cell_6t
Xbit_r59_c192 bl_192 br_192 wl_59 vdd gnd cell_6t
Xbit_r60_c192 bl_192 br_192 wl_60 vdd gnd cell_6t
Xbit_r61_c192 bl_192 br_192 wl_61 vdd gnd cell_6t
Xbit_r62_c192 bl_192 br_192 wl_62 vdd gnd cell_6t
Xbit_r63_c192 bl_192 br_192 wl_63 vdd gnd cell_6t
Xbit_r64_c192 bl_192 br_192 wl_64 vdd gnd cell_6t
Xbit_r65_c192 bl_192 br_192 wl_65 vdd gnd cell_6t
Xbit_r66_c192 bl_192 br_192 wl_66 vdd gnd cell_6t
Xbit_r67_c192 bl_192 br_192 wl_67 vdd gnd cell_6t
Xbit_r68_c192 bl_192 br_192 wl_68 vdd gnd cell_6t
Xbit_r69_c192 bl_192 br_192 wl_69 vdd gnd cell_6t
Xbit_r70_c192 bl_192 br_192 wl_70 vdd gnd cell_6t
Xbit_r71_c192 bl_192 br_192 wl_71 vdd gnd cell_6t
Xbit_r72_c192 bl_192 br_192 wl_72 vdd gnd cell_6t
Xbit_r73_c192 bl_192 br_192 wl_73 vdd gnd cell_6t
Xbit_r74_c192 bl_192 br_192 wl_74 vdd gnd cell_6t
Xbit_r75_c192 bl_192 br_192 wl_75 vdd gnd cell_6t
Xbit_r76_c192 bl_192 br_192 wl_76 vdd gnd cell_6t
Xbit_r77_c192 bl_192 br_192 wl_77 vdd gnd cell_6t
Xbit_r78_c192 bl_192 br_192 wl_78 vdd gnd cell_6t
Xbit_r79_c192 bl_192 br_192 wl_79 vdd gnd cell_6t
Xbit_r80_c192 bl_192 br_192 wl_80 vdd gnd cell_6t
Xbit_r81_c192 bl_192 br_192 wl_81 vdd gnd cell_6t
Xbit_r82_c192 bl_192 br_192 wl_82 vdd gnd cell_6t
Xbit_r83_c192 bl_192 br_192 wl_83 vdd gnd cell_6t
Xbit_r84_c192 bl_192 br_192 wl_84 vdd gnd cell_6t
Xbit_r85_c192 bl_192 br_192 wl_85 vdd gnd cell_6t
Xbit_r86_c192 bl_192 br_192 wl_86 vdd gnd cell_6t
Xbit_r87_c192 bl_192 br_192 wl_87 vdd gnd cell_6t
Xbit_r88_c192 bl_192 br_192 wl_88 vdd gnd cell_6t
Xbit_r89_c192 bl_192 br_192 wl_89 vdd gnd cell_6t
Xbit_r90_c192 bl_192 br_192 wl_90 vdd gnd cell_6t
Xbit_r91_c192 bl_192 br_192 wl_91 vdd gnd cell_6t
Xbit_r92_c192 bl_192 br_192 wl_92 vdd gnd cell_6t
Xbit_r93_c192 bl_192 br_192 wl_93 vdd gnd cell_6t
Xbit_r94_c192 bl_192 br_192 wl_94 vdd gnd cell_6t
Xbit_r95_c192 bl_192 br_192 wl_95 vdd gnd cell_6t
Xbit_r96_c192 bl_192 br_192 wl_96 vdd gnd cell_6t
Xbit_r97_c192 bl_192 br_192 wl_97 vdd gnd cell_6t
Xbit_r98_c192 bl_192 br_192 wl_98 vdd gnd cell_6t
Xbit_r99_c192 bl_192 br_192 wl_99 vdd gnd cell_6t
Xbit_r100_c192 bl_192 br_192 wl_100 vdd gnd cell_6t
Xbit_r101_c192 bl_192 br_192 wl_101 vdd gnd cell_6t
Xbit_r102_c192 bl_192 br_192 wl_102 vdd gnd cell_6t
Xbit_r103_c192 bl_192 br_192 wl_103 vdd gnd cell_6t
Xbit_r104_c192 bl_192 br_192 wl_104 vdd gnd cell_6t
Xbit_r105_c192 bl_192 br_192 wl_105 vdd gnd cell_6t
Xbit_r106_c192 bl_192 br_192 wl_106 vdd gnd cell_6t
Xbit_r107_c192 bl_192 br_192 wl_107 vdd gnd cell_6t
Xbit_r108_c192 bl_192 br_192 wl_108 vdd gnd cell_6t
Xbit_r109_c192 bl_192 br_192 wl_109 vdd gnd cell_6t
Xbit_r110_c192 bl_192 br_192 wl_110 vdd gnd cell_6t
Xbit_r111_c192 bl_192 br_192 wl_111 vdd gnd cell_6t
Xbit_r112_c192 bl_192 br_192 wl_112 vdd gnd cell_6t
Xbit_r113_c192 bl_192 br_192 wl_113 vdd gnd cell_6t
Xbit_r114_c192 bl_192 br_192 wl_114 vdd gnd cell_6t
Xbit_r115_c192 bl_192 br_192 wl_115 vdd gnd cell_6t
Xbit_r116_c192 bl_192 br_192 wl_116 vdd gnd cell_6t
Xbit_r117_c192 bl_192 br_192 wl_117 vdd gnd cell_6t
Xbit_r118_c192 bl_192 br_192 wl_118 vdd gnd cell_6t
Xbit_r119_c192 bl_192 br_192 wl_119 vdd gnd cell_6t
Xbit_r120_c192 bl_192 br_192 wl_120 vdd gnd cell_6t
Xbit_r121_c192 bl_192 br_192 wl_121 vdd gnd cell_6t
Xbit_r122_c192 bl_192 br_192 wl_122 vdd gnd cell_6t
Xbit_r123_c192 bl_192 br_192 wl_123 vdd gnd cell_6t
Xbit_r124_c192 bl_192 br_192 wl_124 vdd gnd cell_6t
Xbit_r125_c192 bl_192 br_192 wl_125 vdd gnd cell_6t
Xbit_r126_c192 bl_192 br_192 wl_126 vdd gnd cell_6t
Xbit_r127_c192 bl_192 br_192 wl_127 vdd gnd cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd cell_6t
Xbit_r1_c193 bl_193 br_193 wl_1 vdd gnd cell_6t
Xbit_r2_c193 bl_193 br_193 wl_2 vdd gnd cell_6t
Xbit_r3_c193 bl_193 br_193 wl_3 vdd gnd cell_6t
Xbit_r4_c193 bl_193 br_193 wl_4 vdd gnd cell_6t
Xbit_r5_c193 bl_193 br_193 wl_5 vdd gnd cell_6t
Xbit_r6_c193 bl_193 br_193 wl_6 vdd gnd cell_6t
Xbit_r7_c193 bl_193 br_193 wl_7 vdd gnd cell_6t
Xbit_r8_c193 bl_193 br_193 wl_8 vdd gnd cell_6t
Xbit_r9_c193 bl_193 br_193 wl_9 vdd gnd cell_6t
Xbit_r10_c193 bl_193 br_193 wl_10 vdd gnd cell_6t
Xbit_r11_c193 bl_193 br_193 wl_11 vdd gnd cell_6t
Xbit_r12_c193 bl_193 br_193 wl_12 vdd gnd cell_6t
Xbit_r13_c193 bl_193 br_193 wl_13 vdd gnd cell_6t
Xbit_r14_c193 bl_193 br_193 wl_14 vdd gnd cell_6t
Xbit_r15_c193 bl_193 br_193 wl_15 vdd gnd cell_6t
Xbit_r16_c193 bl_193 br_193 wl_16 vdd gnd cell_6t
Xbit_r17_c193 bl_193 br_193 wl_17 vdd gnd cell_6t
Xbit_r18_c193 bl_193 br_193 wl_18 vdd gnd cell_6t
Xbit_r19_c193 bl_193 br_193 wl_19 vdd gnd cell_6t
Xbit_r20_c193 bl_193 br_193 wl_20 vdd gnd cell_6t
Xbit_r21_c193 bl_193 br_193 wl_21 vdd gnd cell_6t
Xbit_r22_c193 bl_193 br_193 wl_22 vdd gnd cell_6t
Xbit_r23_c193 bl_193 br_193 wl_23 vdd gnd cell_6t
Xbit_r24_c193 bl_193 br_193 wl_24 vdd gnd cell_6t
Xbit_r25_c193 bl_193 br_193 wl_25 vdd gnd cell_6t
Xbit_r26_c193 bl_193 br_193 wl_26 vdd gnd cell_6t
Xbit_r27_c193 bl_193 br_193 wl_27 vdd gnd cell_6t
Xbit_r28_c193 bl_193 br_193 wl_28 vdd gnd cell_6t
Xbit_r29_c193 bl_193 br_193 wl_29 vdd gnd cell_6t
Xbit_r30_c193 bl_193 br_193 wl_30 vdd gnd cell_6t
Xbit_r31_c193 bl_193 br_193 wl_31 vdd gnd cell_6t
Xbit_r32_c193 bl_193 br_193 wl_32 vdd gnd cell_6t
Xbit_r33_c193 bl_193 br_193 wl_33 vdd gnd cell_6t
Xbit_r34_c193 bl_193 br_193 wl_34 vdd gnd cell_6t
Xbit_r35_c193 bl_193 br_193 wl_35 vdd gnd cell_6t
Xbit_r36_c193 bl_193 br_193 wl_36 vdd gnd cell_6t
Xbit_r37_c193 bl_193 br_193 wl_37 vdd gnd cell_6t
Xbit_r38_c193 bl_193 br_193 wl_38 vdd gnd cell_6t
Xbit_r39_c193 bl_193 br_193 wl_39 vdd gnd cell_6t
Xbit_r40_c193 bl_193 br_193 wl_40 vdd gnd cell_6t
Xbit_r41_c193 bl_193 br_193 wl_41 vdd gnd cell_6t
Xbit_r42_c193 bl_193 br_193 wl_42 vdd gnd cell_6t
Xbit_r43_c193 bl_193 br_193 wl_43 vdd gnd cell_6t
Xbit_r44_c193 bl_193 br_193 wl_44 vdd gnd cell_6t
Xbit_r45_c193 bl_193 br_193 wl_45 vdd gnd cell_6t
Xbit_r46_c193 bl_193 br_193 wl_46 vdd gnd cell_6t
Xbit_r47_c193 bl_193 br_193 wl_47 vdd gnd cell_6t
Xbit_r48_c193 bl_193 br_193 wl_48 vdd gnd cell_6t
Xbit_r49_c193 bl_193 br_193 wl_49 vdd gnd cell_6t
Xbit_r50_c193 bl_193 br_193 wl_50 vdd gnd cell_6t
Xbit_r51_c193 bl_193 br_193 wl_51 vdd gnd cell_6t
Xbit_r52_c193 bl_193 br_193 wl_52 vdd gnd cell_6t
Xbit_r53_c193 bl_193 br_193 wl_53 vdd gnd cell_6t
Xbit_r54_c193 bl_193 br_193 wl_54 vdd gnd cell_6t
Xbit_r55_c193 bl_193 br_193 wl_55 vdd gnd cell_6t
Xbit_r56_c193 bl_193 br_193 wl_56 vdd gnd cell_6t
Xbit_r57_c193 bl_193 br_193 wl_57 vdd gnd cell_6t
Xbit_r58_c193 bl_193 br_193 wl_58 vdd gnd cell_6t
Xbit_r59_c193 bl_193 br_193 wl_59 vdd gnd cell_6t
Xbit_r60_c193 bl_193 br_193 wl_60 vdd gnd cell_6t
Xbit_r61_c193 bl_193 br_193 wl_61 vdd gnd cell_6t
Xbit_r62_c193 bl_193 br_193 wl_62 vdd gnd cell_6t
Xbit_r63_c193 bl_193 br_193 wl_63 vdd gnd cell_6t
Xbit_r64_c193 bl_193 br_193 wl_64 vdd gnd cell_6t
Xbit_r65_c193 bl_193 br_193 wl_65 vdd gnd cell_6t
Xbit_r66_c193 bl_193 br_193 wl_66 vdd gnd cell_6t
Xbit_r67_c193 bl_193 br_193 wl_67 vdd gnd cell_6t
Xbit_r68_c193 bl_193 br_193 wl_68 vdd gnd cell_6t
Xbit_r69_c193 bl_193 br_193 wl_69 vdd gnd cell_6t
Xbit_r70_c193 bl_193 br_193 wl_70 vdd gnd cell_6t
Xbit_r71_c193 bl_193 br_193 wl_71 vdd gnd cell_6t
Xbit_r72_c193 bl_193 br_193 wl_72 vdd gnd cell_6t
Xbit_r73_c193 bl_193 br_193 wl_73 vdd gnd cell_6t
Xbit_r74_c193 bl_193 br_193 wl_74 vdd gnd cell_6t
Xbit_r75_c193 bl_193 br_193 wl_75 vdd gnd cell_6t
Xbit_r76_c193 bl_193 br_193 wl_76 vdd gnd cell_6t
Xbit_r77_c193 bl_193 br_193 wl_77 vdd gnd cell_6t
Xbit_r78_c193 bl_193 br_193 wl_78 vdd gnd cell_6t
Xbit_r79_c193 bl_193 br_193 wl_79 vdd gnd cell_6t
Xbit_r80_c193 bl_193 br_193 wl_80 vdd gnd cell_6t
Xbit_r81_c193 bl_193 br_193 wl_81 vdd gnd cell_6t
Xbit_r82_c193 bl_193 br_193 wl_82 vdd gnd cell_6t
Xbit_r83_c193 bl_193 br_193 wl_83 vdd gnd cell_6t
Xbit_r84_c193 bl_193 br_193 wl_84 vdd gnd cell_6t
Xbit_r85_c193 bl_193 br_193 wl_85 vdd gnd cell_6t
Xbit_r86_c193 bl_193 br_193 wl_86 vdd gnd cell_6t
Xbit_r87_c193 bl_193 br_193 wl_87 vdd gnd cell_6t
Xbit_r88_c193 bl_193 br_193 wl_88 vdd gnd cell_6t
Xbit_r89_c193 bl_193 br_193 wl_89 vdd gnd cell_6t
Xbit_r90_c193 bl_193 br_193 wl_90 vdd gnd cell_6t
Xbit_r91_c193 bl_193 br_193 wl_91 vdd gnd cell_6t
Xbit_r92_c193 bl_193 br_193 wl_92 vdd gnd cell_6t
Xbit_r93_c193 bl_193 br_193 wl_93 vdd gnd cell_6t
Xbit_r94_c193 bl_193 br_193 wl_94 vdd gnd cell_6t
Xbit_r95_c193 bl_193 br_193 wl_95 vdd gnd cell_6t
Xbit_r96_c193 bl_193 br_193 wl_96 vdd gnd cell_6t
Xbit_r97_c193 bl_193 br_193 wl_97 vdd gnd cell_6t
Xbit_r98_c193 bl_193 br_193 wl_98 vdd gnd cell_6t
Xbit_r99_c193 bl_193 br_193 wl_99 vdd gnd cell_6t
Xbit_r100_c193 bl_193 br_193 wl_100 vdd gnd cell_6t
Xbit_r101_c193 bl_193 br_193 wl_101 vdd gnd cell_6t
Xbit_r102_c193 bl_193 br_193 wl_102 vdd gnd cell_6t
Xbit_r103_c193 bl_193 br_193 wl_103 vdd gnd cell_6t
Xbit_r104_c193 bl_193 br_193 wl_104 vdd gnd cell_6t
Xbit_r105_c193 bl_193 br_193 wl_105 vdd gnd cell_6t
Xbit_r106_c193 bl_193 br_193 wl_106 vdd gnd cell_6t
Xbit_r107_c193 bl_193 br_193 wl_107 vdd gnd cell_6t
Xbit_r108_c193 bl_193 br_193 wl_108 vdd gnd cell_6t
Xbit_r109_c193 bl_193 br_193 wl_109 vdd gnd cell_6t
Xbit_r110_c193 bl_193 br_193 wl_110 vdd gnd cell_6t
Xbit_r111_c193 bl_193 br_193 wl_111 vdd gnd cell_6t
Xbit_r112_c193 bl_193 br_193 wl_112 vdd gnd cell_6t
Xbit_r113_c193 bl_193 br_193 wl_113 vdd gnd cell_6t
Xbit_r114_c193 bl_193 br_193 wl_114 vdd gnd cell_6t
Xbit_r115_c193 bl_193 br_193 wl_115 vdd gnd cell_6t
Xbit_r116_c193 bl_193 br_193 wl_116 vdd gnd cell_6t
Xbit_r117_c193 bl_193 br_193 wl_117 vdd gnd cell_6t
Xbit_r118_c193 bl_193 br_193 wl_118 vdd gnd cell_6t
Xbit_r119_c193 bl_193 br_193 wl_119 vdd gnd cell_6t
Xbit_r120_c193 bl_193 br_193 wl_120 vdd gnd cell_6t
Xbit_r121_c193 bl_193 br_193 wl_121 vdd gnd cell_6t
Xbit_r122_c193 bl_193 br_193 wl_122 vdd gnd cell_6t
Xbit_r123_c193 bl_193 br_193 wl_123 vdd gnd cell_6t
Xbit_r124_c193 bl_193 br_193 wl_124 vdd gnd cell_6t
Xbit_r125_c193 bl_193 br_193 wl_125 vdd gnd cell_6t
Xbit_r126_c193 bl_193 br_193 wl_126 vdd gnd cell_6t
Xbit_r127_c193 bl_193 br_193 wl_127 vdd gnd cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd cell_6t
Xbit_r1_c194 bl_194 br_194 wl_1 vdd gnd cell_6t
Xbit_r2_c194 bl_194 br_194 wl_2 vdd gnd cell_6t
Xbit_r3_c194 bl_194 br_194 wl_3 vdd gnd cell_6t
Xbit_r4_c194 bl_194 br_194 wl_4 vdd gnd cell_6t
Xbit_r5_c194 bl_194 br_194 wl_5 vdd gnd cell_6t
Xbit_r6_c194 bl_194 br_194 wl_6 vdd gnd cell_6t
Xbit_r7_c194 bl_194 br_194 wl_7 vdd gnd cell_6t
Xbit_r8_c194 bl_194 br_194 wl_8 vdd gnd cell_6t
Xbit_r9_c194 bl_194 br_194 wl_9 vdd gnd cell_6t
Xbit_r10_c194 bl_194 br_194 wl_10 vdd gnd cell_6t
Xbit_r11_c194 bl_194 br_194 wl_11 vdd gnd cell_6t
Xbit_r12_c194 bl_194 br_194 wl_12 vdd gnd cell_6t
Xbit_r13_c194 bl_194 br_194 wl_13 vdd gnd cell_6t
Xbit_r14_c194 bl_194 br_194 wl_14 vdd gnd cell_6t
Xbit_r15_c194 bl_194 br_194 wl_15 vdd gnd cell_6t
Xbit_r16_c194 bl_194 br_194 wl_16 vdd gnd cell_6t
Xbit_r17_c194 bl_194 br_194 wl_17 vdd gnd cell_6t
Xbit_r18_c194 bl_194 br_194 wl_18 vdd gnd cell_6t
Xbit_r19_c194 bl_194 br_194 wl_19 vdd gnd cell_6t
Xbit_r20_c194 bl_194 br_194 wl_20 vdd gnd cell_6t
Xbit_r21_c194 bl_194 br_194 wl_21 vdd gnd cell_6t
Xbit_r22_c194 bl_194 br_194 wl_22 vdd gnd cell_6t
Xbit_r23_c194 bl_194 br_194 wl_23 vdd gnd cell_6t
Xbit_r24_c194 bl_194 br_194 wl_24 vdd gnd cell_6t
Xbit_r25_c194 bl_194 br_194 wl_25 vdd gnd cell_6t
Xbit_r26_c194 bl_194 br_194 wl_26 vdd gnd cell_6t
Xbit_r27_c194 bl_194 br_194 wl_27 vdd gnd cell_6t
Xbit_r28_c194 bl_194 br_194 wl_28 vdd gnd cell_6t
Xbit_r29_c194 bl_194 br_194 wl_29 vdd gnd cell_6t
Xbit_r30_c194 bl_194 br_194 wl_30 vdd gnd cell_6t
Xbit_r31_c194 bl_194 br_194 wl_31 vdd gnd cell_6t
Xbit_r32_c194 bl_194 br_194 wl_32 vdd gnd cell_6t
Xbit_r33_c194 bl_194 br_194 wl_33 vdd gnd cell_6t
Xbit_r34_c194 bl_194 br_194 wl_34 vdd gnd cell_6t
Xbit_r35_c194 bl_194 br_194 wl_35 vdd gnd cell_6t
Xbit_r36_c194 bl_194 br_194 wl_36 vdd gnd cell_6t
Xbit_r37_c194 bl_194 br_194 wl_37 vdd gnd cell_6t
Xbit_r38_c194 bl_194 br_194 wl_38 vdd gnd cell_6t
Xbit_r39_c194 bl_194 br_194 wl_39 vdd gnd cell_6t
Xbit_r40_c194 bl_194 br_194 wl_40 vdd gnd cell_6t
Xbit_r41_c194 bl_194 br_194 wl_41 vdd gnd cell_6t
Xbit_r42_c194 bl_194 br_194 wl_42 vdd gnd cell_6t
Xbit_r43_c194 bl_194 br_194 wl_43 vdd gnd cell_6t
Xbit_r44_c194 bl_194 br_194 wl_44 vdd gnd cell_6t
Xbit_r45_c194 bl_194 br_194 wl_45 vdd gnd cell_6t
Xbit_r46_c194 bl_194 br_194 wl_46 vdd gnd cell_6t
Xbit_r47_c194 bl_194 br_194 wl_47 vdd gnd cell_6t
Xbit_r48_c194 bl_194 br_194 wl_48 vdd gnd cell_6t
Xbit_r49_c194 bl_194 br_194 wl_49 vdd gnd cell_6t
Xbit_r50_c194 bl_194 br_194 wl_50 vdd gnd cell_6t
Xbit_r51_c194 bl_194 br_194 wl_51 vdd gnd cell_6t
Xbit_r52_c194 bl_194 br_194 wl_52 vdd gnd cell_6t
Xbit_r53_c194 bl_194 br_194 wl_53 vdd gnd cell_6t
Xbit_r54_c194 bl_194 br_194 wl_54 vdd gnd cell_6t
Xbit_r55_c194 bl_194 br_194 wl_55 vdd gnd cell_6t
Xbit_r56_c194 bl_194 br_194 wl_56 vdd gnd cell_6t
Xbit_r57_c194 bl_194 br_194 wl_57 vdd gnd cell_6t
Xbit_r58_c194 bl_194 br_194 wl_58 vdd gnd cell_6t
Xbit_r59_c194 bl_194 br_194 wl_59 vdd gnd cell_6t
Xbit_r60_c194 bl_194 br_194 wl_60 vdd gnd cell_6t
Xbit_r61_c194 bl_194 br_194 wl_61 vdd gnd cell_6t
Xbit_r62_c194 bl_194 br_194 wl_62 vdd gnd cell_6t
Xbit_r63_c194 bl_194 br_194 wl_63 vdd gnd cell_6t
Xbit_r64_c194 bl_194 br_194 wl_64 vdd gnd cell_6t
Xbit_r65_c194 bl_194 br_194 wl_65 vdd gnd cell_6t
Xbit_r66_c194 bl_194 br_194 wl_66 vdd gnd cell_6t
Xbit_r67_c194 bl_194 br_194 wl_67 vdd gnd cell_6t
Xbit_r68_c194 bl_194 br_194 wl_68 vdd gnd cell_6t
Xbit_r69_c194 bl_194 br_194 wl_69 vdd gnd cell_6t
Xbit_r70_c194 bl_194 br_194 wl_70 vdd gnd cell_6t
Xbit_r71_c194 bl_194 br_194 wl_71 vdd gnd cell_6t
Xbit_r72_c194 bl_194 br_194 wl_72 vdd gnd cell_6t
Xbit_r73_c194 bl_194 br_194 wl_73 vdd gnd cell_6t
Xbit_r74_c194 bl_194 br_194 wl_74 vdd gnd cell_6t
Xbit_r75_c194 bl_194 br_194 wl_75 vdd gnd cell_6t
Xbit_r76_c194 bl_194 br_194 wl_76 vdd gnd cell_6t
Xbit_r77_c194 bl_194 br_194 wl_77 vdd gnd cell_6t
Xbit_r78_c194 bl_194 br_194 wl_78 vdd gnd cell_6t
Xbit_r79_c194 bl_194 br_194 wl_79 vdd gnd cell_6t
Xbit_r80_c194 bl_194 br_194 wl_80 vdd gnd cell_6t
Xbit_r81_c194 bl_194 br_194 wl_81 vdd gnd cell_6t
Xbit_r82_c194 bl_194 br_194 wl_82 vdd gnd cell_6t
Xbit_r83_c194 bl_194 br_194 wl_83 vdd gnd cell_6t
Xbit_r84_c194 bl_194 br_194 wl_84 vdd gnd cell_6t
Xbit_r85_c194 bl_194 br_194 wl_85 vdd gnd cell_6t
Xbit_r86_c194 bl_194 br_194 wl_86 vdd gnd cell_6t
Xbit_r87_c194 bl_194 br_194 wl_87 vdd gnd cell_6t
Xbit_r88_c194 bl_194 br_194 wl_88 vdd gnd cell_6t
Xbit_r89_c194 bl_194 br_194 wl_89 vdd gnd cell_6t
Xbit_r90_c194 bl_194 br_194 wl_90 vdd gnd cell_6t
Xbit_r91_c194 bl_194 br_194 wl_91 vdd gnd cell_6t
Xbit_r92_c194 bl_194 br_194 wl_92 vdd gnd cell_6t
Xbit_r93_c194 bl_194 br_194 wl_93 vdd gnd cell_6t
Xbit_r94_c194 bl_194 br_194 wl_94 vdd gnd cell_6t
Xbit_r95_c194 bl_194 br_194 wl_95 vdd gnd cell_6t
Xbit_r96_c194 bl_194 br_194 wl_96 vdd gnd cell_6t
Xbit_r97_c194 bl_194 br_194 wl_97 vdd gnd cell_6t
Xbit_r98_c194 bl_194 br_194 wl_98 vdd gnd cell_6t
Xbit_r99_c194 bl_194 br_194 wl_99 vdd gnd cell_6t
Xbit_r100_c194 bl_194 br_194 wl_100 vdd gnd cell_6t
Xbit_r101_c194 bl_194 br_194 wl_101 vdd gnd cell_6t
Xbit_r102_c194 bl_194 br_194 wl_102 vdd gnd cell_6t
Xbit_r103_c194 bl_194 br_194 wl_103 vdd gnd cell_6t
Xbit_r104_c194 bl_194 br_194 wl_104 vdd gnd cell_6t
Xbit_r105_c194 bl_194 br_194 wl_105 vdd gnd cell_6t
Xbit_r106_c194 bl_194 br_194 wl_106 vdd gnd cell_6t
Xbit_r107_c194 bl_194 br_194 wl_107 vdd gnd cell_6t
Xbit_r108_c194 bl_194 br_194 wl_108 vdd gnd cell_6t
Xbit_r109_c194 bl_194 br_194 wl_109 vdd gnd cell_6t
Xbit_r110_c194 bl_194 br_194 wl_110 vdd gnd cell_6t
Xbit_r111_c194 bl_194 br_194 wl_111 vdd gnd cell_6t
Xbit_r112_c194 bl_194 br_194 wl_112 vdd gnd cell_6t
Xbit_r113_c194 bl_194 br_194 wl_113 vdd gnd cell_6t
Xbit_r114_c194 bl_194 br_194 wl_114 vdd gnd cell_6t
Xbit_r115_c194 bl_194 br_194 wl_115 vdd gnd cell_6t
Xbit_r116_c194 bl_194 br_194 wl_116 vdd gnd cell_6t
Xbit_r117_c194 bl_194 br_194 wl_117 vdd gnd cell_6t
Xbit_r118_c194 bl_194 br_194 wl_118 vdd gnd cell_6t
Xbit_r119_c194 bl_194 br_194 wl_119 vdd gnd cell_6t
Xbit_r120_c194 bl_194 br_194 wl_120 vdd gnd cell_6t
Xbit_r121_c194 bl_194 br_194 wl_121 vdd gnd cell_6t
Xbit_r122_c194 bl_194 br_194 wl_122 vdd gnd cell_6t
Xbit_r123_c194 bl_194 br_194 wl_123 vdd gnd cell_6t
Xbit_r124_c194 bl_194 br_194 wl_124 vdd gnd cell_6t
Xbit_r125_c194 bl_194 br_194 wl_125 vdd gnd cell_6t
Xbit_r126_c194 bl_194 br_194 wl_126 vdd gnd cell_6t
Xbit_r127_c194 bl_194 br_194 wl_127 vdd gnd cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd cell_6t
Xbit_r1_c195 bl_195 br_195 wl_1 vdd gnd cell_6t
Xbit_r2_c195 bl_195 br_195 wl_2 vdd gnd cell_6t
Xbit_r3_c195 bl_195 br_195 wl_3 vdd gnd cell_6t
Xbit_r4_c195 bl_195 br_195 wl_4 vdd gnd cell_6t
Xbit_r5_c195 bl_195 br_195 wl_5 vdd gnd cell_6t
Xbit_r6_c195 bl_195 br_195 wl_6 vdd gnd cell_6t
Xbit_r7_c195 bl_195 br_195 wl_7 vdd gnd cell_6t
Xbit_r8_c195 bl_195 br_195 wl_8 vdd gnd cell_6t
Xbit_r9_c195 bl_195 br_195 wl_9 vdd gnd cell_6t
Xbit_r10_c195 bl_195 br_195 wl_10 vdd gnd cell_6t
Xbit_r11_c195 bl_195 br_195 wl_11 vdd gnd cell_6t
Xbit_r12_c195 bl_195 br_195 wl_12 vdd gnd cell_6t
Xbit_r13_c195 bl_195 br_195 wl_13 vdd gnd cell_6t
Xbit_r14_c195 bl_195 br_195 wl_14 vdd gnd cell_6t
Xbit_r15_c195 bl_195 br_195 wl_15 vdd gnd cell_6t
Xbit_r16_c195 bl_195 br_195 wl_16 vdd gnd cell_6t
Xbit_r17_c195 bl_195 br_195 wl_17 vdd gnd cell_6t
Xbit_r18_c195 bl_195 br_195 wl_18 vdd gnd cell_6t
Xbit_r19_c195 bl_195 br_195 wl_19 vdd gnd cell_6t
Xbit_r20_c195 bl_195 br_195 wl_20 vdd gnd cell_6t
Xbit_r21_c195 bl_195 br_195 wl_21 vdd gnd cell_6t
Xbit_r22_c195 bl_195 br_195 wl_22 vdd gnd cell_6t
Xbit_r23_c195 bl_195 br_195 wl_23 vdd gnd cell_6t
Xbit_r24_c195 bl_195 br_195 wl_24 vdd gnd cell_6t
Xbit_r25_c195 bl_195 br_195 wl_25 vdd gnd cell_6t
Xbit_r26_c195 bl_195 br_195 wl_26 vdd gnd cell_6t
Xbit_r27_c195 bl_195 br_195 wl_27 vdd gnd cell_6t
Xbit_r28_c195 bl_195 br_195 wl_28 vdd gnd cell_6t
Xbit_r29_c195 bl_195 br_195 wl_29 vdd gnd cell_6t
Xbit_r30_c195 bl_195 br_195 wl_30 vdd gnd cell_6t
Xbit_r31_c195 bl_195 br_195 wl_31 vdd gnd cell_6t
Xbit_r32_c195 bl_195 br_195 wl_32 vdd gnd cell_6t
Xbit_r33_c195 bl_195 br_195 wl_33 vdd gnd cell_6t
Xbit_r34_c195 bl_195 br_195 wl_34 vdd gnd cell_6t
Xbit_r35_c195 bl_195 br_195 wl_35 vdd gnd cell_6t
Xbit_r36_c195 bl_195 br_195 wl_36 vdd gnd cell_6t
Xbit_r37_c195 bl_195 br_195 wl_37 vdd gnd cell_6t
Xbit_r38_c195 bl_195 br_195 wl_38 vdd gnd cell_6t
Xbit_r39_c195 bl_195 br_195 wl_39 vdd gnd cell_6t
Xbit_r40_c195 bl_195 br_195 wl_40 vdd gnd cell_6t
Xbit_r41_c195 bl_195 br_195 wl_41 vdd gnd cell_6t
Xbit_r42_c195 bl_195 br_195 wl_42 vdd gnd cell_6t
Xbit_r43_c195 bl_195 br_195 wl_43 vdd gnd cell_6t
Xbit_r44_c195 bl_195 br_195 wl_44 vdd gnd cell_6t
Xbit_r45_c195 bl_195 br_195 wl_45 vdd gnd cell_6t
Xbit_r46_c195 bl_195 br_195 wl_46 vdd gnd cell_6t
Xbit_r47_c195 bl_195 br_195 wl_47 vdd gnd cell_6t
Xbit_r48_c195 bl_195 br_195 wl_48 vdd gnd cell_6t
Xbit_r49_c195 bl_195 br_195 wl_49 vdd gnd cell_6t
Xbit_r50_c195 bl_195 br_195 wl_50 vdd gnd cell_6t
Xbit_r51_c195 bl_195 br_195 wl_51 vdd gnd cell_6t
Xbit_r52_c195 bl_195 br_195 wl_52 vdd gnd cell_6t
Xbit_r53_c195 bl_195 br_195 wl_53 vdd gnd cell_6t
Xbit_r54_c195 bl_195 br_195 wl_54 vdd gnd cell_6t
Xbit_r55_c195 bl_195 br_195 wl_55 vdd gnd cell_6t
Xbit_r56_c195 bl_195 br_195 wl_56 vdd gnd cell_6t
Xbit_r57_c195 bl_195 br_195 wl_57 vdd gnd cell_6t
Xbit_r58_c195 bl_195 br_195 wl_58 vdd gnd cell_6t
Xbit_r59_c195 bl_195 br_195 wl_59 vdd gnd cell_6t
Xbit_r60_c195 bl_195 br_195 wl_60 vdd gnd cell_6t
Xbit_r61_c195 bl_195 br_195 wl_61 vdd gnd cell_6t
Xbit_r62_c195 bl_195 br_195 wl_62 vdd gnd cell_6t
Xbit_r63_c195 bl_195 br_195 wl_63 vdd gnd cell_6t
Xbit_r64_c195 bl_195 br_195 wl_64 vdd gnd cell_6t
Xbit_r65_c195 bl_195 br_195 wl_65 vdd gnd cell_6t
Xbit_r66_c195 bl_195 br_195 wl_66 vdd gnd cell_6t
Xbit_r67_c195 bl_195 br_195 wl_67 vdd gnd cell_6t
Xbit_r68_c195 bl_195 br_195 wl_68 vdd gnd cell_6t
Xbit_r69_c195 bl_195 br_195 wl_69 vdd gnd cell_6t
Xbit_r70_c195 bl_195 br_195 wl_70 vdd gnd cell_6t
Xbit_r71_c195 bl_195 br_195 wl_71 vdd gnd cell_6t
Xbit_r72_c195 bl_195 br_195 wl_72 vdd gnd cell_6t
Xbit_r73_c195 bl_195 br_195 wl_73 vdd gnd cell_6t
Xbit_r74_c195 bl_195 br_195 wl_74 vdd gnd cell_6t
Xbit_r75_c195 bl_195 br_195 wl_75 vdd gnd cell_6t
Xbit_r76_c195 bl_195 br_195 wl_76 vdd gnd cell_6t
Xbit_r77_c195 bl_195 br_195 wl_77 vdd gnd cell_6t
Xbit_r78_c195 bl_195 br_195 wl_78 vdd gnd cell_6t
Xbit_r79_c195 bl_195 br_195 wl_79 vdd gnd cell_6t
Xbit_r80_c195 bl_195 br_195 wl_80 vdd gnd cell_6t
Xbit_r81_c195 bl_195 br_195 wl_81 vdd gnd cell_6t
Xbit_r82_c195 bl_195 br_195 wl_82 vdd gnd cell_6t
Xbit_r83_c195 bl_195 br_195 wl_83 vdd gnd cell_6t
Xbit_r84_c195 bl_195 br_195 wl_84 vdd gnd cell_6t
Xbit_r85_c195 bl_195 br_195 wl_85 vdd gnd cell_6t
Xbit_r86_c195 bl_195 br_195 wl_86 vdd gnd cell_6t
Xbit_r87_c195 bl_195 br_195 wl_87 vdd gnd cell_6t
Xbit_r88_c195 bl_195 br_195 wl_88 vdd gnd cell_6t
Xbit_r89_c195 bl_195 br_195 wl_89 vdd gnd cell_6t
Xbit_r90_c195 bl_195 br_195 wl_90 vdd gnd cell_6t
Xbit_r91_c195 bl_195 br_195 wl_91 vdd gnd cell_6t
Xbit_r92_c195 bl_195 br_195 wl_92 vdd gnd cell_6t
Xbit_r93_c195 bl_195 br_195 wl_93 vdd gnd cell_6t
Xbit_r94_c195 bl_195 br_195 wl_94 vdd gnd cell_6t
Xbit_r95_c195 bl_195 br_195 wl_95 vdd gnd cell_6t
Xbit_r96_c195 bl_195 br_195 wl_96 vdd gnd cell_6t
Xbit_r97_c195 bl_195 br_195 wl_97 vdd gnd cell_6t
Xbit_r98_c195 bl_195 br_195 wl_98 vdd gnd cell_6t
Xbit_r99_c195 bl_195 br_195 wl_99 vdd gnd cell_6t
Xbit_r100_c195 bl_195 br_195 wl_100 vdd gnd cell_6t
Xbit_r101_c195 bl_195 br_195 wl_101 vdd gnd cell_6t
Xbit_r102_c195 bl_195 br_195 wl_102 vdd gnd cell_6t
Xbit_r103_c195 bl_195 br_195 wl_103 vdd gnd cell_6t
Xbit_r104_c195 bl_195 br_195 wl_104 vdd gnd cell_6t
Xbit_r105_c195 bl_195 br_195 wl_105 vdd gnd cell_6t
Xbit_r106_c195 bl_195 br_195 wl_106 vdd gnd cell_6t
Xbit_r107_c195 bl_195 br_195 wl_107 vdd gnd cell_6t
Xbit_r108_c195 bl_195 br_195 wl_108 vdd gnd cell_6t
Xbit_r109_c195 bl_195 br_195 wl_109 vdd gnd cell_6t
Xbit_r110_c195 bl_195 br_195 wl_110 vdd gnd cell_6t
Xbit_r111_c195 bl_195 br_195 wl_111 vdd gnd cell_6t
Xbit_r112_c195 bl_195 br_195 wl_112 vdd gnd cell_6t
Xbit_r113_c195 bl_195 br_195 wl_113 vdd gnd cell_6t
Xbit_r114_c195 bl_195 br_195 wl_114 vdd gnd cell_6t
Xbit_r115_c195 bl_195 br_195 wl_115 vdd gnd cell_6t
Xbit_r116_c195 bl_195 br_195 wl_116 vdd gnd cell_6t
Xbit_r117_c195 bl_195 br_195 wl_117 vdd gnd cell_6t
Xbit_r118_c195 bl_195 br_195 wl_118 vdd gnd cell_6t
Xbit_r119_c195 bl_195 br_195 wl_119 vdd gnd cell_6t
Xbit_r120_c195 bl_195 br_195 wl_120 vdd gnd cell_6t
Xbit_r121_c195 bl_195 br_195 wl_121 vdd gnd cell_6t
Xbit_r122_c195 bl_195 br_195 wl_122 vdd gnd cell_6t
Xbit_r123_c195 bl_195 br_195 wl_123 vdd gnd cell_6t
Xbit_r124_c195 bl_195 br_195 wl_124 vdd gnd cell_6t
Xbit_r125_c195 bl_195 br_195 wl_125 vdd gnd cell_6t
Xbit_r126_c195 bl_195 br_195 wl_126 vdd gnd cell_6t
Xbit_r127_c195 bl_195 br_195 wl_127 vdd gnd cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd cell_6t
Xbit_r1_c196 bl_196 br_196 wl_1 vdd gnd cell_6t
Xbit_r2_c196 bl_196 br_196 wl_2 vdd gnd cell_6t
Xbit_r3_c196 bl_196 br_196 wl_3 vdd gnd cell_6t
Xbit_r4_c196 bl_196 br_196 wl_4 vdd gnd cell_6t
Xbit_r5_c196 bl_196 br_196 wl_5 vdd gnd cell_6t
Xbit_r6_c196 bl_196 br_196 wl_6 vdd gnd cell_6t
Xbit_r7_c196 bl_196 br_196 wl_7 vdd gnd cell_6t
Xbit_r8_c196 bl_196 br_196 wl_8 vdd gnd cell_6t
Xbit_r9_c196 bl_196 br_196 wl_9 vdd gnd cell_6t
Xbit_r10_c196 bl_196 br_196 wl_10 vdd gnd cell_6t
Xbit_r11_c196 bl_196 br_196 wl_11 vdd gnd cell_6t
Xbit_r12_c196 bl_196 br_196 wl_12 vdd gnd cell_6t
Xbit_r13_c196 bl_196 br_196 wl_13 vdd gnd cell_6t
Xbit_r14_c196 bl_196 br_196 wl_14 vdd gnd cell_6t
Xbit_r15_c196 bl_196 br_196 wl_15 vdd gnd cell_6t
Xbit_r16_c196 bl_196 br_196 wl_16 vdd gnd cell_6t
Xbit_r17_c196 bl_196 br_196 wl_17 vdd gnd cell_6t
Xbit_r18_c196 bl_196 br_196 wl_18 vdd gnd cell_6t
Xbit_r19_c196 bl_196 br_196 wl_19 vdd gnd cell_6t
Xbit_r20_c196 bl_196 br_196 wl_20 vdd gnd cell_6t
Xbit_r21_c196 bl_196 br_196 wl_21 vdd gnd cell_6t
Xbit_r22_c196 bl_196 br_196 wl_22 vdd gnd cell_6t
Xbit_r23_c196 bl_196 br_196 wl_23 vdd gnd cell_6t
Xbit_r24_c196 bl_196 br_196 wl_24 vdd gnd cell_6t
Xbit_r25_c196 bl_196 br_196 wl_25 vdd gnd cell_6t
Xbit_r26_c196 bl_196 br_196 wl_26 vdd gnd cell_6t
Xbit_r27_c196 bl_196 br_196 wl_27 vdd gnd cell_6t
Xbit_r28_c196 bl_196 br_196 wl_28 vdd gnd cell_6t
Xbit_r29_c196 bl_196 br_196 wl_29 vdd gnd cell_6t
Xbit_r30_c196 bl_196 br_196 wl_30 vdd gnd cell_6t
Xbit_r31_c196 bl_196 br_196 wl_31 vdd gnd cell_6t
Xbit_r32_c196 bl_196 br_196 wl_32 vdd gnd cell_6t
Xbit_r33_c196 bl_196 br_196 wl_33 vdd gnd cell_6t
Xbit_r34_c196 bl_196 br_196 wl_34 vdd gnd cell_6t
Xbit_r35_c196 bl_196 br_196 wl_35 vdd gnd cell_6t
Xbit_r36_c196 bl_196 br_196 wl_36 vdd gnd cell_6t
Xbit_r37_c196 bl_196 br_196 wl_37 vdd gnd cell_6t
Xbit_r38_c196 bl_196 br_196 wl_38 vdd gnd cell_6t
Xbit_r39_c196 bl_196 br_196 wl_39 vdd gnd cell_6t
Xbit_r40_c196 bl_196 br_196 wl_40 vdd gnd cell_6t
Xbit_r41_c196 bl_196 br_196 wl_41 vdd gnd cell_6t
Xbit_r42_c196 bl_196 br_196 wl_42 vdd gnd cell_6t
Xbit_r43_c196 bl_196 br_196 wl_43 vdd gnd cell_6t
Xbit_r44_c196 bl_196 br_196 wl_44 vdd gnd cell_6t
Xbit_r45_c196 bl_196 br_196 wl_45 vdd gnd cell_6t
Xbit_r46_c196 bl_196 br_196 wl_46 vdd gnd cell_6t
Xbit_r47_c196 bl_196 br_196 wl_47 vdd gnd cell_6t
Xbit_r48_c196 bl_196 br_196 wl_48 vdd gnd cell_6t
Xbit_r49_c196 bl_196 br_196 wl_49 vdd gnd cell_6t
Xbit_r50_c196 bl_196 br_196 wl_50 vdd gnd cell_6t
Xbit_r51_c196 bl_196 br_196 wl_51 vdd gnd cell_6t
Xbit_r52_c196 bl_196 br_196 wl_52 vdd gnd cell_6t
Xbit_r53_c196 bl_196 br_196 wl_53 vdd gnd cell_6t
Xbit_r54_c196 bl_196 br_196 wl_54 vdd gnd cell_6t
Xbit_r55_c196 bl_196 br_196 wl_55 vdd gnd cell_6t
Xbit_r56_c196 bl_196 br_196 wl_56 vdd gnd cell_6t
Xbit_r57_c196 bl_196 br_196 wl_57 vdd gnd cell_6t
Xbit_r58_c196 bl_196 br_196 wl_58 vdd gnd cell_6t
Xbit_r59_c196 bl_196 br_196 wl_59 vdd gnd cell_6t
Xbit_r60_c196 bl_196 br_196 wl_60 vdd gnd cell_6t
Xbit_r61_c196 bl_196 br_196 wl_61 vdd gnd cell_6t
Xbit_r62_c196 bl_196 br_196 wl_62 vdd gnd cell_6t
Xbit_r63_c196 bl_196 br_196 wl_63 vdd gnd cell_6t
Xbit_r64_c196 bl_196 br_196 wl_64 vdd gnd cell_6t
Xbit_r65_c196 bl_196 br_196 wl_65 vdd gnd cell_6t
Xbit_r66_c196 bl_196 br_196 wl_66 vdd gnd cell_6t
Xbit_r67_c196 bl_196 br_196 wl_67 vdd gnd cell_6t
Xbit_r68_c196 bl_196 br_196 wl_68 vdd gnd cell_6t
Xbit_r69_c196 bl_196 br_196 wl_69 vdd gnd cell_6t
Xbit_r70_c196 bl_196 br_196 wl_70 vdd gnd cell_6t
Xbit_r71_c196 bl_196 br_196 wl_71 vdd gnd cell_6t
Xbit_r72_c196 bl_196 br_196 wl_72 vdd gnd cell_6t
Xbit_r73_c196 bl_196 br_196 wl_73 vdd gnd cell_6t
Xbit_r74_c196 bl_196 br_196 wl_74 vdd gnd cell_6t
Xbit_r75_c196 bl_196 br_196 wl_75 vdd gnd cell_6t
Xbit_r76_c196 bl_196 br_196 wl_76 vdd gnd cell_6t
Xbit_r77_c196 bl_196 br_196 wl_77 vdd gnd cell_6t
Xbit_r78_c196 bl_196 br_196 wl_78 vdd gnd cell_6t
Xbit_r79_c196 bl_196 br_196 wl_79 vdd gnd cell_6t
Xbit_r80_c196 bl_196 br_196 wl_80 vdd gnd cell_6t
Xbit_r81_c196 bl_196 br_196 wl_81 vdd gnd cell_6t
Xbit_r82_c196 bl_196 br_196 wl_82 vdd gnd cell_6t
Xbit_r83_c196 bl_196 br_196 wl_83 vdd gnd cell_6t
Xbit_r84_c196 bl_196 br_196 wl_84 vdd gnd cell_6t
Xbit_r85_c196 bl_196 br_196 wl_85 vdd gnd cell_6t
Xbit_r86_c196 bl_196 br_196 wl_86 vdd gnd cell_6t
Xbit_r87_c196 bl_196 br_196 wl_87 vdd gnd cell_6t
Xbit_r88_c196 bl_196 br_196 wl_88 vdd gnd cell_6t
Xbit_r89_c196 bl_196 br_196 wl_89 vdd gnd cell_6t
Xbit_r90_c196 bl_196 br_196 wl_90 vdd gnd cell_6t
Xbit_r91_c196 bl_196 br_196 wl_91 vdd gnd cell_6t
Xbit_r92_c196 bl_196 br_196 wl_92 vdd gnd cell_6t
Xbit_r93_c196 bl_196 br_196 wl_93 vdd gnd cell_6t
Xbit_r94_c196 bl_196 br_196 wl_94 vdd gnd cell_6t
Xbit_r95_c196 bl_196 br_196 wl_95 vdd gnd cell_6t
Xbit_r96_c196 bl_196 br_196 wl_96 vdd gnd cell_6t
Xbit_r97_c196 bl_196 br_196 wl_97 vdd gnd cell_6t
Xbit_r98_c196 bl_196 br_196 wl_98 vdd gnd cell_6t
Xbit_r99_c196 bl_196 br_196 wl_99 vdd gnd cell_6t
Xbit_r100_c196 bl_196 br_196 wl_100 vdd gnd cell_6t
Xbit_r101_c196 bl_196 br_196 wl_101 vdd gnd cell_6t
Xbit_r102_c196 bl_196 br_196 wl_102 vdd gnd cell_6t
Xbit_r103_c196 bl_196 br_196 wl_103 vdd gnd cell_6t
Xbit_r104_c196 bl_196 br_196 wl_104 vdd gnd cell_6t
Xbit_r105_c196 bl_196 br_196 wl_105 vdd gnd cell_6t
Xbit_r106_c196 bl_196 br_196 wl_106 vdd gnd cell_6t
Xbit_r107_c196 bl_196 br_196 wl_107 vdd gnd cell_6t
Xbit_r108_c196 bl_196 br_196 wl_108 vdd gnd cell_6t
Xbit_r109_c196 bl_196 br_196 wl_109 vdd gnd cell_6t
Xbit_r110_c196 bl_196 br_196 wl_110 vdd gnd cell_6t
Xbit_r111_c196 bl_196 br_196 wl_111 vdd gnd cell_6t
Xbit_r112_c196 bl_196 br_196 wl_112 vdd gnd cell_6t
Xbit_r113_c196 bl_196 br_196 wl_113 vdd gnd cell_6t
Xbit_r114_c196 bl_196 br_196 wl_114 vdd gnd cell_6t
Xbit_r115_c196 bl_196 br_196 wl_115 vdd gnd cell_6t
Xbit_r116_c196 bl_196 br_196 wl_116 vdd gnd cell_6t
Xbit_r117_c196 bl_196 br_196 wl_117 vdd gnd cell_6t
Xbit_r118_c196 bl_196 br_196 wl_118 vdd gnd cell_6t
Xbit_r119_c196 bl_196 br_196 wl_119 vdd gnd cell_6t
Xbit_r120_c196 bl_196 br_196 wl_120 vdd gnd cell_6t
Xbit_r121_c196 bl_196 br_196 wl_121 vdd gnd cell_6t
Xbit_r122_c196 bl_196 br_196 wl_122 vdd gnd cell_6t
Xbit_r123_c196 bl_196 br_196 wl_123 vdd gnd cell_6t
Xbit_r124_c196 bl_196 br_196 wl_124 vdd gnd cell_6t
Xbit_r125_c196 bl_196 br_196 wl_125 vdd gnd cell_6t
Xbit_r126_c196 bl_196 br_196 wl_126 vdd gnd cell_6t
Xbit_r127_c196 bl_196 br_196 wl_127 vdd gnd cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd cell_6t
Xbit_r1_c197 bl_197 br_197 wl_1 vdd gnd cell_6t
Xbit_r2_c197 bl_197 br_197 wl_2 vdd gnd cell_6t
Xbit_r3_c197 bl_197 br_197 wl_3 vdd gnd cell_6t
Xbit_r4_c197 bl_197 br_197 wl_4 vdd gnd cell_6t
Xbit_r5_c197 bl_197 br_197 wl_5 vdd gnd cell_6t
Xbit_r6_c197 bl_197 br_197 wl_6 vdd gnd cell_6t
Xbit_r7_c197 bl_197 br_197 wl_7 vdd gnd cell_6t
Xbit_r8_c197 bl_197 br_197 wl_8 vdd gnd cell_6t
Xbit_r9_c197 bl_197 br_197 wl_9 vdd gnd cell_6t
Xbit_r10_c197 bl_197 br_197 wl_10 vdd gnd cell_6t
Xbit_r11_c197 bl_197 br_197 wl_11 vdd gnd cell_6t
Xbit_r12_c197 bl_197 br_197 wl_12 vdd gnd cell_6t
Xbit_r13_c197 bl_197 br_197 wl_13 vdd gnd cell_6t
Xbit_r14_c197 bl_197 br_197 wl_14 vdd gnd cell_6t
Xbit_r15_c197 bl_197 br_197 wl_15 vdd gnd cell_6t
Xbit_r16_c197 bl_197 br_197 wl_16 vdd gnd cell_6t
Xbit_r17_c197 bl_197 br_197 wl_17 vdd gnd cell_6t
Xbit_r18_c197 bl_197 br_197 wl_18 vdd gnd cell_6t
Xbit_r19_c197 bl_197 br_197 wl_19 vdd gnd cell_6t
Xbit_r20_c197 bl_197 br_197 wl_20 vdd gnd cell_6t
Xbit_r21_c197 bl_197 br_197 wl_21 vdd gnd cell_6t
Xbit_r22_c197 bl_197 br_197 wl_22 vdd gnd cell_6t
Xbit_r23_c197 bl_197 br_197 wl_23 vdd gnd cell_6t
Xbit_r24_c197 bl_197 br_197 wl_24 vdd gnd cell_6t
Xbit_r25_c197 bl_197 br_197 wl_25 vdd gnd cell_6t
Xbit_r26_c197 bl_197 br_197 wl_26 vdd gnd cell_6t
Xbit_r27_c197 bl_197 br_197 wl_27 vdd gnd cell_6t
Xbit_r28_c197 bl_197 br_197 wl_28 vdd gnd cell_6t
Xbit_r29_c197 bl_197 br_197 wl_29 vdd gnd cell_6t
Xbit_r30_c197 bl_197 br_197 wl_30 vdd gnd cell_6t
Xbit_r31_c197 bl_197 br_197 wl_31 vdd gnd cell_6t
Xbit_r32_c197 bl_197 br_197 wl_32 vdd gnd cell_6t
Xbit_r33_c197 bl_197 br_197 wl_33 vdd gnd cell_6t
Xbit_r34_c197 bl_197 br_197 wl_34 vdd gnd cell_6t
Xbit_r35_c197 bl_197 br_197 wl_35 vdd gnd cell_6t
Xbit_r36_c197 bl_197 br_197 wl_36 vdd gnd cell_6t
Xbit_r37_c197 bl_197 br_197 wl_37 vdd gnd cell_6t
Xbit_r38_c197 bl_197 br_197 wl_38 vdd gnd cell_6t
Xbit_r39_c197 bl_197 br_197 wl_39 vdd gnd cell_6t
Xbit_r40_c197 bl_197 br_197 wl_40 vdd gnd cell_6t
Xbit_r41_c197 bl_197 br_197 wl_41 vdd gnd cell_6t
Xbit_r42_c197 bl_197 br_197 wl_42 vdd gnd cell_6t
Xbit_r43_c197 bl_197 br_197 wl_43 vdd gnd cell_6t
Xbit_r44_c197 bl_197 br_197 wl_44 vdd gnd cell_6t
Xbit_r45_c197 bl_197 br_197 wl_45 vdd gnd cell_6t
Xbit_r46_c197 bl_197 br_197 wl_46 vdd gnd cell_6t
Xbit_r47_c197 bl_197 br_197 wl_47 vdd gnd cell_6t
Xbit_r48_c197 bl_197 br_197 wl_48 vdd gnd cell_6t
Xbit_r49_c197 bl_197 br_197 wl_49 vdd gnd cell_6t
Xbit_r50_c197 bl_197 br_197 wl_50 vdd gnd cell_6t
Xbit_r51_c197 bl_197 br_197 wl_51 vdd gnd cell_6t
Xbit_r52_c197 bl_197 br_197 wl_52 vdd gnd cell_6t
Xbit_r53_c197 bl_197 br_197 wl_53 vdd gnd cell_6t
Xbit_r54_c197 bl_197 br_197 wl_54 vdd gnd cell_6t
Xbit_r55_c197 bl_197 br_197 wl_55 vdd gnd cell_6t
Xbit_r56_c197 bl_197 br_197 wl_56 vdd gnd cell_6t
Xbit_r57_c197 bl_197 br_197 wl_57 vdd gnd cell_6t
Xbit_r58_c197 bl_197 br_197 wl_58 vdd gnd cell_6t
Xbit_r59_c197 bl_197 br_197 wl_59 vdd gnd cell_6t
Xbit_r60_c197 bl_197 br_197 wl_60 vdd gnd cell_6t
Xbit_r61_c197 bl_197 br_197 wl_61 vdd gnd cell_6t
Xbit_r62_c197 bl_197 br_197 wl_62 vdd gnd cell_6t
Xbit_r63_c197 bl_197 br_197 wl_63 vdd gnd cell_6t
Xbit_r64_c197 bl_197 br_197 wl_64 vdd gnd cell_6t
Xbit_r65_c197 bl_197 br_197 wl_65 vdd gnd cell_6t
Xbit_r66_c197 bl_197 br_197 wl_66 vdd gnd cell_6t
Xbit_r67_c197 bl_197 br_197 wl_67 vdd gnd cell_6t
Xbit_r68_c197 bl_197 br_197 wl_68 vdd gnd cell_6t
Xbit_r69_c197 bl_197 br_197 wl_69 vdd gnd cell_6t
Xbit_r70_c197 bl_197 br_197 wl_70 vdd gnd cell_6t
Xbit_r71_c197 bl_197 br_197 wl_71 vdd gnd cell_6t
Xbit_r72_c197 bl_197 br_197 wl_72 vdd gnd cell_6t
Xbit_r73_c197 bl_197 br_197 wl_73 vdd gnd cell_6t
Xbit_r74_c197 bl_197 br_197 wl_74 vdd gnd cell_6t
Xbit_r75_c197 bl_197 br_197 wl_75 vdd gnd cell_6t
Xbit_r76_c197 bl_197 br_197 wl_76 vdd gnd cell_6t
Xbit_r77_c197 bl_197 br_197 wl_77 vdd gnd cell_6t
Xbit_r78_c197 bl_197 br_197 wl_78 vdd gnd cell_6t
Xbit_r79_c197 bl_197 br_197 wl_79 vdd gnd cell_6t
Xbit_r80_c197 bl_197 br_197 wl_80 vdd gnd cell_6t
Xbit_r81_c197 bl_197 br_197 wl_81 vdd gnd cell_6t
Xbit_r82_c197 bl_197 br_197 wl_82 vdd gnd cell_6t
Xbit_r83_c197 bl_197 br_197 wl_83 vdd gnd cell_6t
Xbit_r84_c197 bl_197 br_197 wl_84 vdd gnd cell_6t
Xbit_r85_c197 bl_197 br_197 wl_85 vdd gnd cell_6t
Xbit_r86_c197 bl_197 br_197 wl_86 vdd gnd cell_6t
Xbit_r87_c197 bl_197 br_197 wl_87 vdd gnd cell_6t
Xbit_r88_c197 bl_197 br_197 wl_88 vdd gnd cell_6t
Xbit_r89_c197 bl_197 br_197 wl_89 vdd gnd cell_6t
Xbit_r90_c197 bl_197 br_197 wl_90 vdd gnd cell_6t
Xbit_r91_c197 bl_197 br_197 wl_91 vdd gnd cell_6t
Xbit_r92_c197 bl_197 br_197 wl_92 vdd gnd cell_6t
Xbit_r93_c197 bl_197 br_197 wl_93 vdd gnd cell_6t
Xbit_r94_c197 bl_197 br_197 wl_94 vdd gnd cell_6t
Xbit_r95_c197 bl_197 br_197 wl_95 vdd gnd cell_6t
Xbit_r96_c197 bl_197 br_197 wl_96 vdd gnd cell_6t
Xbit_r97_c197 bl_197 br_197 wl_97 vdd gnd cell_6t
Xbit_r98_c197 bl_197 br_197 wl_98 vdd gnd cell_6t
Xbit_r99_c197 bl_197 br_197 wl_99 vdd gnd cell_6t
Xbit_r100_c197 bl_197 br_197 wl_100 vdd gnd cell_6t
Xbit_r101_c197 bl_197 br_197 wl_101 vdd gnd cell_6t
Xbit_r102_c197 bl_197 br_197 wl_102 vdd gnd cell_6t
Xbit_r103_c197 bl_197 br_197 wl_103 vdd gnd cell_6t
Xbit_r104_c197 bl_197 br_197 wl_104 vdd gnd cell_6t
Xbit_r105_c197 bl_197 br_197 wl_105 vdd gnd cell_6t
Xbit_r106_c197 bl_197 br_197 wl_106 vdd gnd cell_6t
Xbit_r107_c197 bl_197 br_197 wl_107 vdd gnd cell_6t
Xbit_r108_c197 bl_197 br_197 wl_108 vdd gnd cell_6t
Xbit_r109_c197 bl_197 br_197 wl_109 vdd gnd cell_6t
Xbit_r110_c197 bl_197 br_197 wl_110 vdd gnd cell_6t
Xbit_r111_c197 bl_197 br_197 wl_111 vdd gnd cell_6t
Xbit_r112_c197 bl_197 br_197 wl_112 vdd gnd cell_6t
Xbit_r113_c197 bl_197 br_197 wl_113 vdd gnd cell_6t
Xbit_r114_c197 bl_197 br_197 wl_114 vdd gnd cell_6t
Xbit_r115_c197 bl_197 br_197 wl_115 vdd gnd cell_6t
Xbit_r116_c197 bl_197 br_197 wl_116 vdd gnd cell_6t
Xbit_r117_c197 bl_197 br_197 wl_117 vdd gnd cell_6t
Xbit_r118_c197 bl_197 br_197 wl_118 vdd gnd cell_6t
Xbit_r119_c197 bl_197 br_197 wl_119 vdd gnd cell_6t
Xbit_r120_c197 bl_197 br_197 wl_120 vdd gnd cell_6t
Xbit_r121_c197 bl_197 br_197 wl_121 vdd gnd cell_6t
Xbit_r122_c197 bl_197 br_197 wl_122 vdd gnd cell_6t
Xbit_r123_c197 bl_197 br_197 wl_123 vdd gnd cell_6t
Xbit_r124_c197 bl_197 br_197 wl_124 vdd gnd cell_6t
Xbit_r125_c197 bl_197 br_197 wl_125 vdd gnd cell_6t
Xbit_r126_c197 bl_197 br_197 wl_126 vdd gnd cell_6t
Xbit_r127_c197 bl_197 br_197 wl_127 vdd gnd cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd cell_6t
Xbit_r1_c198 bl_198 br_198 wl_1 vdd gnd cell_6t
Xbit_r2_c198 bl_198 br_198 wl_2 vdd gnd cell_6t
Xbit_r3_c198 bl_198 br_198 wl_3 vdd gnd cell_6t
Xbit_r4_c198 bl_198 br_198 wl_4 vdd gnd cell_6t
Xbit_r5_c198 bl_198 br_198 wl_5 vdd gnd cell_6t
Xbit_r6_c198 bl_198 br_198 wl_6 vdd gnd cell_6t
Xbit_r7_c198 bl_198 br_198 wl_7 vdd gnd cell_6t
Xbit_r8_c198 bl_198 br_198 wl_8 vdd gnd cell_6t
Xbit_r9_c198 bl_198 br_198 wl_9 vdd gnd cell_6t
Xbit_r10_c198 bl_198 br_198 wl_10 vdd gnd cell_6t
Xbit_r11_c198 bl_198 br_198 wl_11 vdd gnd cell_6t
Xbit_r12_c198 bl_198 br_198 wl_12 vdd gnd cell_6t
Xbit_r13_c198 bl_198 br_198 wl_13 vdd gnd cell_6t
Xbit_r14_c198 bl_198 br_198 wl_14 vdd gnd cell_6t
Xbit_r15_c198 bl_198 br_198 wl_15 vdd gnd cell_6t
Xbit_r16_c198 bl_198 br_198 wl_16 vdd gnd cell_6t
Xbit_r17_c198 bl_198 br_198 wl_17 vdd gnd cell_6t
Xbit_r18_c198 bl_198 br_198 wl_18 vdd gnd cell_6t
Xbit_r19_c198 bl_198 br_198 wl_19 vdd gnd cell_6t
Xbit_r20_c198 bl_198 br_198 wl_20 vdd gnd cell_6t
Xbit_r21_c198 bl_198 br_198 wl_21 vdd gnd cell_6t
Xbit_r22_c198 bl_198 br_198 wl_22 vdd gnd cell_6t
Xbit_r23_c198 bl_198 br_198 wl_23 vdd gnd cell_6t
Xbit_r24_c198 bl_198 br_198 wl_24 vdd gnd cell_6t
Xbit_r25_c198 bl_198 br_198 wl_25 vdd gnd cell_6t
Xbit_r26_c198 bl_198 br_198 wl_26 vdd gnd cell_6t
Xbit_r27_c198 bl_198 br_198 wl_27 vdd gnd cell_6t
Xbit_r28_c198 bl_198 br_198 wl_28 vdd gnd cell_6t
Xbit_r29_c198 bl_198 br_198 wl_29 vdd gnd cell_6t
Xbit_r30_c198 bl_198 br_198 wl_30 vdd gnd cell_6t
Xbit_r31_c198 bl_198 br_198 wl_31 vdd gnd cell_6t
Xbit_r32_c198 bl_198 br_198 wl_32 vdd gnd cell_6t
Xbit_r33_c198 bl_198 br_198 wl_33 vdd gnd cell_6t
Xbit_r34_c198 bl_198 br_198 wl_34 vdd gnd cell_6t
Xbit_r35_c198 bl_198 br_198 wl_35 vdd gnd cell_6t
Xbit_r36_c198 bl_198 br_198 wl_36 vdd gnd cell_6t
Xbit_r37_c198 bl_198 br_198 wl_37 vdd gnd cell_6t
Xbit_r38_c198 bl_198 br_198 wl_38 vdd gnd cell_6t
Xbit_r39_c198 bl_198 br_198 wl_39 vdd gnd cell_6t
Xbit_r40_c198 bl_198 br_198 wl_40 vdd gnd cell_6t
Xbit_r41_c198 bl_198 br_198 wl_41 vdd gnd cell_6t
Xbit_r42_c198 bl_198 br_198 wl_42 vdd gnd cell_6t
Xbit_r43_c198 bl_198 br_198 wl_43 vdd gnd cell_6t
Xbit_r44_c198 bl_198 br_198 wl_44 vdd gnd cell_6t
Xbit_r45_c198 bl_198 br_198 wl_45 vdd gnd cell_6t
Xbit_r46_c198 bl_198 br_198 wl_46 vdd gnd cell_6t
Xbit_r47_c198 bl_198 br_198 wl_47 vdd gnd cell_6t
Xbit_r48_c198 bl_198 br_198 wl_48 vdd gnd cell_6t
Xbit_r49_c198 bl_198 br_198 wl_49 vdd gnd cell_6t
Xbit_r50_c198 bl_198 br_198 wl_50 vdd gnd cell_6t
Xbit_r51_c198 bl_198 br_198 wl_51 vdd gnd cell_6t
Xbit_r52_c198 bl_198 br_198 wl_52 vdd gnd cell_6t
Xbit_r53_c198 bl_198 br_198 wl_53 vdd gnd cell_6t
Xbit_r54_c198 bl_198 br_198 wl_54 vdd gnd cell_6t
Xbit_r55_c198 bl_198 br_198 wl_55 vdd gnd cell_6t
Xbit_r56_c198 bl_198 br_198 wl_56 vdd gnd cell_6t
Xbit_r57_c198 bl_198 br_198 wl_57 vdd gnd cell_6t
Xbit_r58_c198 bl_198 br_198 wl_58 vdd gnd cell_6t
Xbit_r59_c198 bl_198 br_198 wl_59 vdd gnd cell_6t
Xbit_r60_c198 bl_198 br_198 wl_60 vdd gnd cell_6t
Xbit_r61_c198 bl_198 br_198 wl_61 vdd gnd cell_6t
Xbit_r62_c198 bl_198 br_198 wl_62 vdd gnd cell_6t
Xbit_r63_c198 bl_198 br_198 wl_63 vdd gnd cell_6t
Xbit_r64_c198 bl_198 br_198 wl_64 vdd gnd cell_6t
Xbit_r65_c198 bl_198 br_198 wl_65 vdd gnd cell_6t
Xbit_r66_c198 bl_198 br_198 wl_66 vdd gnd cell_6t
Xbit_r67_c198 bl_198 br_198 wl_67 vdd gnd cell_6t
Xbit_r68_c198 bl_198 br_198 wl_68 vdd gnd cell_6t
Xbit_r69_c198 bl_198 br_198 wl_69 vdd gnd cell_6t
Xbit_r70_c198 bl_198 br_198 wl_70 vdd gnd cell_6t
Xbit_r71_c198 bl_198 br_198 wl_71 vdd gnd cell_6t
Xbit_r72_c198 bl_198 br_198 wl_72 vdd gnd cell_6t
Xbit_r73_c198 bl_198 br_198 wl_73 vdd gnd cell_6t
Xbit_r74_c198 bl_198 br_198 wl_74 vdd gnd cell_6t
Xbit_r75_c198 bl_198 br_198 wl_75 vdd gnd cell_6t
Xbit_r76_c198 bl_198 br_198 wl_76 vdd gnd cell_6t
Xbit_r77_c198 bl_198 br_198 wl_77 vdd gnd cell_6t
Xbit_r78_c198 bl_198 br_198 wl_78 vdd gnd cell_6t
Xbit_r79_c198 bl_198 br_198 wl_79 vdd gnd cell_6t
Xbit_r80_c198 bl_198 br_198 wl_80 vdd gnd cell_6t
Xbit_r81_c198 bl_198 br_198 wl_81 vdd gnd cell_6t
Xbit_r82_c198 bl_198 br_198 wl_82 vdd gnd cell_6t
Xbit_r83_c198 bl_198 br_198 wl_83 vdd gnd cell_6t
Xbit_r84_c198 bl_198 br_198 wl_84 vdd gnd cell_6t
Xbit_r85_c198 bl_198 br_198 wl_85 vdd gnd cell_6t
Xbit_r86_c198 bl_198 br_198 wl_86 vdd gnd cell_6t
Xbit_r87_c198 bl_198 br_198 wl_87 vdd gnd cell_6t
Xbit_r88_c198 bl_198 br_198 wl_88 vdd gnd cell_6t
Xbit_r89_c198 bl_198 br_198 wl_89 vdd gnd cell_6t
Xbit_r90_c198 bl_198 br_198 wl_90 vdd gnd cell_6t
Xbit_r91_c198 bl_198 br_198 wl_91 vdd gnd cell_6t
Xbit_r92_c198 bl_198 br_198 wl_92 vdd gnd cell_6t
Xbit_r93_c198 bl_198 br_198 wl_93 vdd gnd cell_6t
Xbit_r94_c198 bl_198 br_198 wl_94 vdd gnd cell_6t
Xbit_r95_c198 bl_198 br_198 wl_95 vdd gnd cell_6t
Xbit_r96_c198 bl_198 br_198 wl_96 vdd gnd cell_6t
Xbit_r97_c198 bl_198 br_198 wl_97 vdd gnd cell_6t
Xbit_r98_c198 bl_198 br_198 wl_98 vdd gnd cell_6t
Xbit_r99_c198 bl_198 br_198 wl_99 vdd gnd cell_6t
Xbit_r100_c198 bl_198 br_198 wl_100 vdd gnd cell_6t
Xbit_r101_c198 bl_198 br_198 wl_101 vdd gnd cell_6t
Xbit_r102_c198 bl_198 br_198 wl_102 vdd gnd cell_6t
Xbit_r103_c198 bl_198 br_198 wl_103 vdd gnd cell_6t
Xbit_r104_c198 bl_198 br_198 wl_104 vdd gnd cell_6t
Xbit_r105_c198 bl_198 br_198 wl_105 vdd gnd cell_6t
Xbit_r106_c198 bl_198 br_198 wl_106 vdd gnd cell_6t
Xbit_r107_c198 bl_198 br_198 wl_107 vdd gnd cell_6t
Xbit_r108_c198 bl_198 br_198 wl_108 vdd gnd cell_6t
Xbit_r109_c198 bl_198 br_198 wl_109 vdd gnd cell_6t
Xbit_r110_c198 bl_198 br_198 wl_110 vdd gnd cell_6t
Xbit_r111_c198 bl_198 br_198 wl_111 vdd gnd cell_6t
Xbit_r112_c198 bl_198 br_198 wl_112 vdd gnd cell_6t
Xbit_r113_c198 bl_198 br_198 wl_113 vdd gnd cell_6t
Xbit_r114_c198 bl_198 br_198 wl_114 vdd gnd cell_6t
Xbit_r115_c198 bl_198 br_198 wl_115 vdd gnd cell_6t
Xbit_r116_c198 bl_198 br_198 wl_116 vdd gnd cell_6t
Xbit_r117_c198 bl_198 br_198 wl_117 vdd gnd cell_6t
Xbit_r118_c198 bl_198 br_198 wl_118 vdd gnd cell_6t
Xbit_r119_c198 bl_198 br_198 wl_119 vdd gnd cell_6t
Xbit_r120_c198 bl_198 br_198 wl_120 vdd gnd cell_6t
Xbit_r121_c198 bl_198 br_198 wl_121 vdd gnd cell_6t
Xbit_r122_c198 bl_198 br_198 wl_122 vdd gnd cell_6t
Xbit_r123_c198 bl_198 br_198 wl_123 vdd gnd cell_6t
Xbit_r124_c198 bl_198 br_198 wl_124 vdd gnd cell_6t
Xbit_r125_c198 bl_198 br_198 wl_125 vdd gnd cell_6t
Xbit_r126_c198 bl_198 br_198 wl_126 vdd gnd cell_6t
Xbit_r127_c198 bl_198 br_198 wl_127 vdd gnd cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd cell_6t
Xbit_r1_c199 bl_199 br_199 wl_1 vdd gnd cell_6t
Xbit_r2_c199 bl_199 br_199 wl_2 vdd gnd cell_6t
Xbit_r3_c199 bl_199 br_199 wl_3 vdd gnd cell_6t
Xbit_r4_c199 bl_199 br_199 wl_4 vdd gnd cell_6t
Xbit_r5_c199 bl_199 br_199 wl_5 vdd gnd cell_6t
Xbit_r6_c199 bl_199 br_199 wl_6 vdd gnd cell_6t
Xbit_r7_c199 bl_199 br_199 wl_7 vdd gnd cell_6t
Xbit_r8_c199 bl_199 br_199 wl_8 vdd gnd cell_6t
Xbit_r9_c199 bl_199 br_199 wl_9 vdd gnd cell_6t
Xbit_r10_c199 bl_199 br_199 wl_10 vdd gnd cell_6t
Xbit_r11_c199 bl_199 br_199 wl_11 vdd gnd cell_6t
Xbit_r12_c199 bl_199 br_199 wl_12 vdd gnd cell_6t
Xbit_r13_c199 bl_199 br_199 wl_13 vdd gnd cell_6t
Xbit_r14_c199 bl_199 br_199 wl_14 vdd gnd cell_6t
Xbit_r15_c199 bl_199 br_199 wl_15 vdd gnd cell_6t
Xbit_r16_c199 bl_199 br_199 wl_16 vdd gnd cell_6t
Xbit_r17_c199 bl_199 br_199 wl_17 vdd gnd cell_6t
Xbit_r18_c199 bl_199 br_199 wl_18 vdd gnd cell_6t
Xbit_r19_c199 bl_199 br_199 wl_19 vdd gnd cell_6t
Xbit_r20_c199 bl_199 br_199 wl_20 vdd gnd cell_6t
Xbit_r21_c199 bl_199 br_199 wl_21 vdd gnd cell_6t
Xbit_r22_c199 bl_199 br_199 wl_22 vdd gnd cell_6t
Xbit_r23_c199 bl_199 br_199 wl_23 vdd gnd cell_6t
Xbit_r24_c199 bl_199 br_199 wl_24 vdd gnd cell_6t
Xbit_r25_c199 bl_199 br_199 wl_25 vdd gnd cell_6t
Xbit_r26_c199 bl_199 br_199 wl_26 vdd gnd cell_6t
Xbit_r27_c199 bl_199 br_199 wl_27 vdd gnd cell_6t
Xbit_r28_c199 bl_199 br_199 wl_28 vdd gnd cell_6t
Xbit_r29_c199 bl_199 br_199 wl_29 vdd gnd cell_6t
Xbit_r30_c199 bl_199 br_199 wl_30 vdd gnd cell_6t
Xbit_r31_c199 bl_199 br_199 wl_31 vdd gnd cell_6t
Xbit_r32_c199 bl_199 br_199 wl_32 vdd gnd cell_6t
Xbit_r33_c199 bl_199 br_199 wl_33 vdd gnd cell_6t
Xbit_r34_c199 bl_199 br_199 wl_34 vdd gnd cell_6t
Xbit_r35_c199 bl_199 br_199 wl_35 vdd gnd cell_6t
Xbit_r36_c199 bl_199 br_199 wl_36 vdd gnd cell_6t
Xbit_r37_c199 bl_199 br_199 wl_37 vdd gnd cell_6t
Xbit_r38_c199 bl_199 br_199 wl_38 vdd gnd cell_6t
Xbit_r39_c199 bl_199 br_199 wl_39 vdd gnd cell_6t
Xbit_r40_c199 bl_199 br_199 wl_40 vdd gnd cell_6t
Xbit_r41_c199 bl_199 br_199 wl_41 vdd gnd cell_6t
Xbit_r42_c199 bl_199 br_199 wl_42 vdd gnd cell_6t
Xbit_r43_c199 bl_199 br_199 wl_43 vdd gnd cell_6t
Xbit_r44_c199 bl_199 br_199 wl_44 vdd gnd cell_6t
Xbit_r45_c199 bl_199 br_199 wl_45 vdd gnd cell_6t
Xbit_r46_c199 bl_199 br_199 wl_46 vdd gnd cell_6t
Xbit_r47_c199 bl_199 br_199 wl_47 vdd gnd cell_6t
Xbit_r48_c199 bl_199 br_199 wl_48 vdd gnd cell_6t
Xbit_r49_c199 bl_199 br_199 wl_49 vdd gnd cell_6t
Xbit_r50_c199 bl_199 br_199 wl_50 vdd gnd cell_6t
Xbit_r51_c199 bl_199 br_199 wl_51 vdd gnd cell_6t
Xbit_r52_c199 bl_199 br_199 wl_52 vdd gnd cell_6t
Xbit_r53_c199 bl_199 br_199 wl_53 vdd gnd cell_6t
Xbit_r54_c199 bl_199 br_199 wl_54 vdd gnd cell_6t
Xbit_r55_c199 bl_199 br_199 wl_55 vdd gnd cell_6t
Xbit_r56_c199 bl_199 br_199 wl_56 vdd gnd cell_6t
Xbit_r57_c199 bl_199 br_199 wl_57 vdd gnd cell_6t
Xbit_r58_c199 bl_199 br_199 wl_58 vdd gnd cell_6t
Xbit_r59_c199 bl_199 br_199 wl_59 vdd gnd cell_6t
Xbit_r60_c199 bl_199 br_199 wl_60 vdd gnd cell_6t
Xbit_r61_c199 bl_199 br_199 wl_61 vdd gnd cell_6t
Xbit_r62_c199 bl_199 br_199 wl_62 vdd gnd cell_6t
Xbit_r63_c199 bl_199 br_199 wl_63 vdd gnd cell_6t
Xbit_r64_c199 bl_199 br_199 wl_64 vdd gnd cell_6t
Xbit_r65_c199 bl_199 br_199 wl_65 vdd gnd cell_6t
Xbit_r66_c199 bl_199 br_199 wl_66 vdd gnd cell_6t
Xbit_r67_c199 bl_199 br_199 wl_67 vdd gnd cell_6t
Xbit_r68_c199 bl_199 br_199 wl_68 vdd gnd cell_6t
Xbit_r69_c199 bl_199 br_199 wl_69 vdd gnd cell_6t
Xbit_r70_c199 bl_199 br_199 wl_70 vdd gnd cell_6t
Xbit_r71_c199 bl_199 br_199 wl_71 vdd gnd cell_6t
Xbit_r72_c199 bl_199 br_199 wl_72 vdd gnd cell_6t
Xbit_r73_c199 bl_199 br_199 wl_73 vdd gnd cell_6t
Xbit_r74_c199 bl_199 br_199 wl_74 vdd gnd cell_6t
Xbit_r75_c199 bl_199 br_199 wl_75 vdd gnd cell_6t
Xbit_r76_c199 bl_199 br_199 wl_76 vdd gnd cell_6t
Xbit_r77_c199 bl_199 br_199 wl_77 vdd gnd cell_6t
Xbit_r78_c199 bl_199 br_199 wl_78 vdd gnd cell_6t
Xbit_r79_c199 bl_199 br_199 wl_79 vdd gnd cell_6t
Xbit_r80_c199 bl_199 br_199 wl_80 vdd gnd cell_6t
Xbit_r81_c199 bl_199 br_199 wl_81 vdd gnd cell_6t
Xbit_r82_c199 bl_199 br_199 wl_82 vdd gnd cell_6t
Xbit_r83_c199 bl_199 br_199 wl_83 vdd gnd cell_6t
Xbit_r84_c199 bl_199 br_199 wl_84 vdd gnd cell_6t
Xbit_r85_c199 bl_199 br_199 wl_85 vdd gnd cell_6t
Xbit_r86_c199 bl_199 br_199 wl_86 vdd gnd cell_6t
Xbit_r87_c199 bl_199 br_199 wl_87 vdd gnd cell_6t
Xbit_r88_c199 bl_199 br_199 wl_88 vdd gnd cell_6t
Xbit_r89_c199 bl_199 br_199 wl_89 vdd gnd cell_6t
Xbit_r90_c199 bl_199 br_199 wl_90 vdd gnd cell_6t
Xbit_r91_c199 bl_199 br_199 wl_91 vdd gnd cell_6t
Xbit_r92_c199 bl_199 br_199 wl_92 vdd gnd cell_6t
Xbit_r93_c199 bl_199 br_199 wl_93 vdd gnd cell_6t
Xbit_r94_c199 bl_199 br_199 wl_94 vdd gnd cell_6t
Xbit_r95_c199 bl_199 br_199 wl_95 vdd gnd cell_6t
Xbit_r96_c199 bl_199 br_199 wl_96 vdd gnd cell_6t
Xbit_r97_c199 bl_199 br_199 wl_97 vdd gnd cell_6t
Xbit_r98_c199 bl_199 br_199 wl_98 vdd gnd cell_6t
Xbit_r99_c199 bl_199 br_199 wl_99 vdd gnd cell_6t
Xbit_r100_c199 bl_199 br_199 wl_100 vdd gnd cell_6t
Xbit_r101_c199 bl_199 br_199 wl_101 vdd gnd cell_6t
Xbit_r102_c199 bl_199 br_199 wl_102 vdd gnd cell_6t
Xbit_r103_c199 bl_199 br_199 wl_103 vdd gnd cell_6t
Xbit_r104_c199 bl_199 br_199 wl_104 vdd gnd cell_6t
Xbit_r105_c199 bl_199 br_199 wl_105 vdd gnd cell_6t
Xbit_r106_c199 bl_199 br_199 wl_106 vdd gnd cell_6t
Xbit_r107_c199 bl_199 br_199 wl_107 vdd gnd cell_6t
Xbit_r108_c199 bl_199 br_199 wl_108 vdd gnd cell_6t
Xbit_r109_c199 bl_199 br_199 wl_109 vdd gnd cell_6t
Xbit_r110_c199 bl_199 br_199 wl_110 vdd gnd cell_6t
Xbit_r111_c199 bl_199 br_199 wl_111 vdd gnd cell_6t
Xbit_r112_c199 bl_199 br_199 wl_112 vdd gnd cell_6t
Xbit_r113_c199 bl_199 br_199 wl_113 vdd gnd cell_6t
Xbit_r114_c199 bl_199 br_199 wl_114 vdd gnd cell_6t
Xbit_r115_c199 bl_199 br_199 wl_115 vdd gnd cell_6t
Xbit_r116_c199 bl_199 br_199 wl_116 vdd gnd cell_6t
Xbit_r117_c199 bl_199 br_199 wl_117 vdd gnd cell_6t
Xbit_r118_c199 bl_199 br_199 wl_118 vdd gnd cell_6t
Xbit_r119_c199 bl_199 br_199 wl_119 vdd gnd cell_6t
Xbit_r120_c199 bl_199 br_199 wl_120 vdd gnd cell_6t
Xbit_r121_c199 bl_199 br_199 wl_121 vdd gnd cell_6t
Xbit_r122_c199 bl_199 br_199 wl_122 vdd gnd cell_6t
Xbit_r123_c199 bl_199 br_199 wl_123 vdd gnd cell_6t
Xbit_r124_c199 bl_199 br_199 wl_124 vdd gnd cell_6t
Xbit_r125_c199 bl_199 br_199 wl_125 vdd gnd cell_6t
Xbit_r126_c199 bl_199 br_199 wl_126 vdd gnd cell_6t
Xbit_r127_c199 bl_199 br_199 wl_127 vdd gnd cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd cell_6t
Xbit_r1_c200 bl_200 br_200 wl_1 vdd gnd cell_6t
Xbit_r2_c200 bl_200 br_200 wl_2 vdd gnd cell_6t
Xbit_r3_c200 bl_200 br_200 wl_3 vdd gnd cell_6t
Xbit_r4_c200 bl_200 br_200 wl_4 vdd gnd cell_6t
Xbit_r5_c200 bl_200 br_200 wl_5 vdd gnd cell_6t
Xbit_r6_c200 bl_200 br_200 wl_6 vdd gnd cell_6t
Xbit_r7_c200 bl_200 br_200 wl_7 vdd gnd cell_6t
Xbit_r8_c200 bl_200 br_200 wl_8 vdd gnd cell_6t
Xbit_r9_c200 bl_200 br_200 wl_9 vdd gnd cell_6t
Xbit_r10_c200 bl_200 br_200 wl_10 vdd gnd cell_6t
Xbit_r11_c200 bl_200 br_200 wl_11 vdd gnd cell_6t
Xbit_r12_c200 bl_200 br_200 wl_12 vdd gnd cell_6t
Xbit_r13_c200 bl_200 br_200 wl_13 vdd gnd cell_6t
Xbit_r14_c200 bl_200 br_200 wl_14 vdd gnd cell_6t
Xbit_r15_c200 bl_200 br_200 wl_15 vdd gnd cell_6t
Xbit_r16_c200 bl_200 br_200 wl_16 vdd gnd cell_6t
Xbit_r17_c200 bl_200 br_200 wl_17 vdd gnd cell_6t
Xbit_r18_c200 bl_200 br_200 wl_18 vdd gnd cell_6t
Xbit_r19_c200 bl_200 br_200 wl_19 vdd gnd cell_6t
Xbit_r20_c200 bl_200 br_200 wl_20 vdd gnd cell_6t
Xbit_r21_c200 bl_200 br_200 wl_21 vdd gnd cell_6t
Xbit_r22_c200 bl_200 br_200 wl_22 vdd gnd cell_6t
Xbit_r23_c200 bl_200 br_200 wl_23 vdd gnd cell_6t
Xbit_r24_c200 bl_200 br_200 wl_24 vdd gnd cell_6t
Xbit_r25_c200 bl_200 br_200 wl_25 vdd gnd cell_6t
Xbit_r26_c200 bl_200 br_200 wl_26 vdd gnd cell_6t
Xbit_r27_c200 bl_200 br_200 wl_27 vdd gnd cell_6t
Xbit_r28_c200 bl_200 br_200 wl_28 vdd gnd cell_6t
Xbit_r29_c200 bl_200 br_200 wl_29 vdd gnd cell_6t
Xbit_r30_c200 bl_200 br_200 wl_30 vdd gnd cell_6t
Xbit_r31_c200 bl_200 br_200 wl_31 vdd gnd cell_6t
Xbit_r32_c200 bl_200 br_200 wl_32 vdd gnd cell_6t
Xbit_r33_c200 bl_200 br_200 wl_33 vdd gnd cell_6t
Xbit_r34_c200 bl_200 br_200 wl_34 vdd gnd cell_6t
Xbit_r35_c200 bl_200 br_200 wl_35 vdd gnd cell_6t
Xbit_r36_c200 bl_200 br_200 wl_36 vdd gnd cell_6t
Xbit_r37_c200 bl_200 br_200 wl_37 vdd gnd cell_6t
Xbit_r38_c200 bl_200 br_200 wl_38 vdd gnd cell_6t
Xbit_r39_c200 bl_200 br_200 wl_39 vdd gnd cell_6t
Xbit_r40_c200 bl_200 br_200 wl_40 vdd gnd cell_6t
Xbit_r41_c200 bl_200 br_200 wl_41 vdd gnd cell_6t
Xbit_r42_c200 bl_200 br_200 wl_42 vdd gnd cell_6t
Xbit_r43_c200 bl_200 br_200 wl_43 vdd gnd cell_6t
Xbit_r44_c200 bl_200 br_200 wl_44 vdd gnd cell_6t
Xbit_r45_c200 bl_200 br_200 wl_45 vdd gnd cell_6t
Xbit_r46_c200 bl_200 br_200 wl_46 vdd gnd cell_6t
Xbit_r47_c200 bl_200 br_200 wl_47 vdd gnd cell_6t
Xbit_r48_c200 bl_200 br_200 wl_48 vdd gnd cell_6t
Xbit_r49_c200 bl_200 br_200 wl_49 vdd gnd cell_6t
Xbit_r50_c200 bl_200 br_200 wl_50 vdd gnd cell_6t
Xbit_r51_c200 bl_200 br_200 wl_51 vdd gnd cell_6t
Xbit_r52_c200 bl_200 br_200 wl_52 vdd gnd cell_6t
Xbit_r53_c200 bl_200 br_200 wl_53 vdd gnd cell_6t
Xbit_r54_c200 bl_200 br_200 wl_54 vdd gnd cell_6t
Xbit_r55_c200 bl_200 br_200 wl_55 vdd gnd cell_6t
Xbit_r56_c200 bl_200 br_200 wl_56 vdd gnd cell_6t
Xbit_r57_c200 bl_200 br_200 wl_57 vdd gnd cell_6t
Xbit_r58_c200 bl_200 br_200 wl_58 vdd gnd cell_6t
Xbit_r59_c200 bl_200 br_200 wl_59 vdd gnd cell_6t
Xbit_r60_c200 bl_200 br_200 wl_60 vdd gnd cell_6t
Xbit_r61_c200 bl_200 br_200 wl_61 vdd gnd cell_6t
Xbit_r62_c200 bl_200 br_200 wl_62 vdd gnd cell_6t
Xbit_r63_c200 bl_200 br_200 wl_63 vdd gnd cell_6t
Xbit_r64_c200 bl_200 br_200 wl_64 vdd gnd cell_6t
Xbit_r65_c200 bl_200 br_200 wl_65 vdd gnd cell_6t
Xbit_r66_c200 bl_200 br_200 wl_66 vdd gnd cell_6t
Xbit_r67_c200 bl_200 br_200 wl_67 vdd gnd cell_6t
Xbit_r68_c200 bl_200 br_200 wl_68 vdd gnd cell_6t
Xbit_r69_c200 bl_200 br_200 wl_69 vdd gnd cell_6t
Xbit_r70_c200 bl_200 br_200 wl_70 vdd gnd cell_6t
Xbit_r71_c200 bl_200 br_200 wl_71 vdd gnd cell_6t
Xbit_r72_c200 bl_200 br_200 wl_72 vdd gnd cell_6t
Xbit_r73_c200 bl_200 br_200 wl_73 vdd gnd cell_6t
Xbit_r74_c200 bl_200 br_200 wl_74 vdd gnd cell_6t
Xbit_r75_c200 bl_200 br_200 wl_75 vdd gnd cell_6t
Xbit_r76_c200 bl_200 br_200 wl_76 vdd gnd cell_6t
Xbit_r77_c200 bl_200 br_200 wl_77 vdd gnd cell_6t
Xbit_r78_c200 bl_200 br_200 wl_78 vdd gnd cell_6t
Xbit_r79_c200 bl_200 br_200 wl_79 vdd gnd cell_6t
Xbit_r80_c200 bl_200 br_200 wl_80 vdd gnd cell_6t
Xbit_r81_c200 bl_200 br_200 wl_81 vdd gnd cell_6t
Xbit_r82_c200 bl_200 br_200 wl_82 vdd gnd cell_6t
Xbit_r83_c200 bl_200 br_200 wl_83 vdd gnd cell_6t
Xbit_r84_c200 bl_200 br_200 wl_84 vdd gnd cell_6t
Xbit_r85_c200 bl_200 br_200 wl_85 vdd gnd cell_6t
Xbit_r86_c200 bl_200 br_200 wl_86 vdd gnd cell_6t
Xbit_r87_c200 bl_200 br_200 wl_87 vdd gnd cell_6t
Xbit_r88_c200 bl_200 br_200 wl_88 vdd gnd cell_6t
Xbit_r89_c200 bl_200 br_200 wl_89 vdd gnd cell_6t
Xbit_r90_c200 bl_200 br_200 wl_90 vdd gnd cell_6t
Xbit_r91_c200 bl_200 br_200 wl_91 vdd gnd cell_6t
Xbit_r92_c200 bl_200 br_200 wl_92 vdd gnd cell_6t
Xbit_r93_c200 bl_200 br_200 wl_93 vdd gnd cell_6t
Xbit_r94_c200 bl_200 br_200 wl_94 vdd gnd cell_6t
Xbit_r95_c200 bl_200 br_200 wl_95 vdd gnd cell_6t
Xbit_r96_c200 bl_200 br_200 wl_96 vdd gnd cell_6t
Xbit_r97_c200 bl_200 br_200 wl_97 vdd gnd cell_6t
Xbit_r98_c200 bl_200 br_200 wl_98 vdd gnd cell_6t
Xbit_r99_c200 bl_200 br_200 wl_99 vdd gnd cell_6t
Xbit_r100_c200 bl_200 br_200 wl_100 vdd gnd cell_6t
Xbit_r101_c200 bl_200 br_200 wl_101 vdd gnd cell_6t
Xbit_r102_c200 bl_200 br_200 wl_102 vdd gnd cell_6t
Xbit_r103_c200 bl_200 br_200 wl_103 vdd gnd cell_6t
Xbit_r104_c200 bl_200 br_200 wl_104 vdd gnd cell_6t
Xbit_r105_c200 bl_200 br_200 wl_105 vdd gnd cell_6t
Xbit_r106_c200 bl_200 br_200 wl_106 vdd gnd cell_6t
Xbit_r107_c200 bl_200 br_200 wl_107 vdd gnd cell_6t
Xbit_r108_c200 bl_200 br_200 wl_108 vdd gnd cell_6t
Xbit_r109_c200 bl_200 br_200 wl_109 vdd gnd cell_6t
Xbit_r110_c200 bl_200 br_200 wl_110 vdd gnd cell_6t
Xbit_r111_c200 bl_200 br_200 wl_111 vdd gnd cell_6t
Xbit_r112_c200 bl_200 br_200 wl_112 vdd gnd cell_6t
Xbit_r113_c200 bl_200 br_200 wl_113 vdd gnd cell_6t
Xbit_r114_c200 bl_200 br_200 wl_114 vdd gnd cell_6t
Xbit_r115_c200 bl_200 br_200 wl_115 vdd gnd cell_6t
Xbit_r116_c200 bl_200 br_200 wl_116 vdd gnd cell_6t
Xbit_r117_c200 bl_200 br_200 wl_117 vdd gnd cell_6t
Xbit_r118_c200 bl_200 br_200 wl_118 vdd gnd cell_6t
Xbit_r119_c200 bl_200 br_200 wl_119 vdd gnd cell_6t
Xbit_r120_c200 bl_200 br_200 wl_120 vdd gnd cell_6t
Xbit_r121_c200 bl_200 br_200 wl_121 vdd gnd cell_6t
Xbit_r122_c200 bl_200 br_200 wl_122 vdd gnd cell_6t
Xbit_r123_c200 bl_200 br_200 wl_123 vdd gnd cell_6t
Xbit_r124_c200 bl_200 br_200 wl_124 vdd gnd cell_6t
Xbit_r125_c200 bl_200 br_200 wl_125 vdd gnd cell_6t
Xbit_r126_c200 bl_200 br_200 wl_126 vdd gnd cell_6t
Xbit_r127_c200 bl_200 br_200 wl_127 vdd gnd cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd cell_6t
Xbit_r1_c201 bl_201 br_201 wl_1 vdd gnd cell_6t
Xbit_r2_c201 bl_201 br_201 wl_2 vdd gnd cell_6t
Xbit_r3_c201 bl_201 br_201 wl_3 vdd gnd cell_6t
Xbit_r4_c201 bl_201 br_201 wl_4 vdd gnd cell_6t
Xbit_r5_c201 bl_201 br_201 wl_5 vdd gnd cell_6t
Xbit_r6_c201 bl_201 br_201 wl_6 vdd gnd cell_6t
Xbit_r7_c201 bl_201 br_201 wl_7 vdd gnd cell_6t
Xbit_r8_c201 bl_201 br_201 wl_8 vdd gnd cell_6t
Xbit_r9_c201 bl_201 br_201 wl_9 vdd gnd cell_6t
Xbit_r10_c201 bl_201 br_201 wl_10 vdd gnd cell_6t
Xbit_r11_c201 bl_201 br_201 wl_11 vdd gnd cell_6t
Xbit_r12_c201 bl_201 br_201 wl_12 vdd gnd cell_6t
Xbit_r13_c201 bl_201 br_201 wl_13 vdd gnd cell_6t
Xbit_r14_c201 bl_201 br_201 wl_14 vdd gnd cell_6t
Xbit_r15_c201 bl_201 br_201 wl_15 vdd gnd cell_6t
Xbit_r16_c201 bl_201 br_201 wl_16 vdd gnd cell_6t
Xbit_r17_c201 bl_201 br_201 wl_17 vdd gnd cell_6t
Xbit_r18_c201 bl_201 br_201 wl_18 vdd gnd cell_6t
Xbit_r19_c201 bl_201 br_201 wl_19 vdd gnd cell_6t
Xbit_r20_c201 bl_201 br_201 wl_20 vdd gnd cell_6t
Xbit_r21_c201 bl_201 br_201 wl_21 vdd gnd cell_6t
Xbit_r22_c201 bl_201 br_201 wl_22 vdd gnd cell_6t
Xbit_r23_c201 bl_201 br_201 wl_23 vdd gnd cell_6t
Xbit_r24_c201 bl_201 br_201 wl_24 vdd gnd cell_6t
Xbit_r25_c201 bl_201 br_201 wl_25 vdd gnd cell_6t
Xbit_r26_c201 bl_201 br_201 wl_26 vdd gnd cell_6t
Xbit_r27_c201 bl_201 br_201 wl_27 vdd gnd cell_6t
Xbit_r28_c201 bl_201 br_201 wl_28 vdd gnd cell_6t
Xbit_r29_c201 bl_201 br_201 wl_29 vdd gnd cell_6t
Xbit_r30_c201 bl_201 br_201 wl_30 vdd gnd cell_6t
Xbit_r31_c201 bl_201 br_201 wl_31 vdd gnd cell_6t
Xbit_r32_c201 bl_201 br_201 wl_32 vdd gnd cell_6t
Xbit_r33_c201 bl_201 br_201 wl_33 vdd gnd cell_6t
Xbit_r34_c201 bl_201 br_201 wl_34 vdd gnd cell_6t
Xbit_r35_c201 bl_201 br_201 wl_35 vdd gnd cell_6t
Xbit_r36_c201 bl_201 br_201 wl_36 vdd gnd cell_6t
Xbit_r37_c201 bl_201 br_201 wl_37 vdd gnd cell_6t
Xbit_r38_c201 bl_201 br_201 wl_38 vdd gnd cell_6t
Xbit_r39_c201 bl_201 br_201 wl_39 vdd gnd cell_6t
Xbit_r40_c201 bl_201 br_201 wl_40 vdd gnd cell_6t
Xbit_r41_c201 bl_201 br_201 wl_41 vdd gnd cell_6t
Xbit_r42_c201 bl_201 br_201 wl_42 vdd gnd cell_6t
Xbit_r43_c201 bl_201 br_201 wl_43 vdd gnd cell_6t
Xbit_r44_c201 bl_201 br_201 wl_44 vdd gnd cell_6t
Xbit_r45_c201 bl_201 br_201 wl_45 vdd gnd cell_6t
Xbit_r46_c201 bl_201 br_201 wl_46 vdd gnd cell_6t
Xbit_r47_c201 bl_201 br_201 wl_47 vdd gnd cell_6t
Xbit_r48_c201 bl_201 br_201 wl_48 vdd gnd cell_6t
Xbit_r49_c201 bl_201 br_201 wl_49 vdd gnd cell_6t
Xbit_r50_c201 bl_201 br_201 wl_50 vdd gnd cell_6t
Xbit_r51_c201 bl_201 br_201 wl_51 vdd gnd cell_6t
Xbit_r52_c201 bl_201 br_201 wl_52 vdd gnd cell_6t
Xbit_r53_c201 bl_201 br_201 wl_53 vdd gnd cell_6t
Xbit_r54_c201 bl_201 br_201 wl_54 vdd gnd cell_6t
Xbit_r55_c201 bl_201 br_201 wl_55 vdd gnd cell_6t
Xbit_r56_c201 bl_201 br_201 wl_56 vdd gnd cell_6t
Xbit_r57_c201 bl_201 br_201 wl_57 vdd gnd cell_6t
Xbit_r58_c201 bl_201 br_201 wl_58 vdd gnd cell_6t
Xbit_r59_c201 bl_201 br_201 wl_59 vdd gnd cell_6t
Xbit_r60_c201 bl_201 br_201 wl_60 vdd gnd cell_6t
Xbit_r61_c201 bl_201 br_201 wl_61 vdd gnd cell_6t
Xbit_r62_c201 bl_201 br_201 wl_62 vdd gnd cell_6t
Xbit_r63_c201 bl_201 br_201 wl_63 vdd gnd cell_6t
Xbit_r64_c201 bl_201 br_201 wl_64 vdd gnd cell_6t
Xbit_r65_c201 bl_201 br_201 wl_65 vdd gnd cell_6t
Xbit_r66_c201 bl_201 br_201 wl_66 vdd gnd cell_6t
Xbit_r67_c201 bl_201 br_201 wl_67 vdd gnd cell_6t
Xbit_r68_c201 bl_201 br_201 wl_68 vdd gnd cell_6t
Xbit_r69_c201 bl_201 br_201 wl_69 vdd gnd cell_6t
Xbit_r70_c201 bl_201 br_201 wl_70 vdd gnd cell_6t
Xbit_r71_c201 bl_201 br_201 wl_71 vdd gnd cell_6t
Xbit_r72_c201 bl_201 br_201 wl_72 vdd gnd cell_6t
Xbit_r73_c201 bl_201 br_201 wl_73 vdd gnd cell_6t
Xbit_r74_c201 bl_201 br_201 wl_74 vdd gnd cell_6t
Xbit_r75_c201 bl_201 br_201 wl_75 vdd gnd cell_6t
Xbit_r76_c201 bl_201 br_201 wl_76 vdd gnd cell_6t
Xbit_r77_c201 bl_201 br_201 wl_77 vdd gnd cell_6t
Xbit_r78_c201 bl_201 br_201 wl_78 vdd gnd cell_6t
Xbit_r79_c201 bl_201 br_201 wl_79 vdd gnd cell_6t
Xbit_r80_c201 bl_201 br_201 wl_80 vdd gnd cell_6t
Xbit_r81_c201 bl_201 br_201 wl_81 vdd gnd cell_6t
Xbit_r82_c201 bl_201 br_201 wl_82 vdd gnd cell_6t
Xbit_r83_c201 bl_201 br_201 wl_83 vdd gnd cell_6t
Xbit_r84_c201 bl_201 br_201 wl_84 vdd gnd cell_6t
Xbit_r85_c201 bl_201 br_201 wl_85 vdd gnd cell_6t
Xbit_r86_c201 bl_201 br_201 wl_86 vdd gnd cell_6t
Xbit_r87_c201 bl_201 br_201 wl_87 vdd gnd cell_6t
Xbit_r88_c201 bl_201 br_201 wl_88 vdd gnd cell_6t
Xbit_r89_c201 bl_201 br_201 wl_89 vdd gnd cell_6t
Xbit_r90_c201 bl_201 br_201 wl_90 vdd gnd cell_6t
Xbit_r91_c201 bl_201 br_201 wl_91 vdd gnd cell_6t
Xbit_r92_c201 bl_201 br_201 wl_92 vdd gnd cell_6t
Xbit_r93_c201 bl_201 br_201 wl_93 vdd gnd cell_6t
Xbit_r94_c201 bl_201 br_201 wl_94 vdd gnd cell_6t
Xbit_r95_c201 bl_201 br_201 wl_95 vdd gnd cell_6t
Xbit_r96_c201 bl_201 br_201 wl_96 vdd gnd cell_6t
Xbit_r97_c201 bl_201 br_201 wl_97 vdd gnd cell_6t
Xbit_r98_c201 bl_201 br_201 wl_98 vdd gnd cell_6t
Xbit_r99_c201 bl_201 br_201 wl_99 vdd gnd cell_6t
Xbit_r100_c201 bl_201 br_201 wl_100 vdd gnd cell_6t
Xbit_r101_c201 bl_201 br_201 wl_101 vdd gnd cell_6t
Xbit_r102_c201 bl_201 br_201 wl_102 vdd gnd cell_6t
Xbit_r103_c201 bl_201 br_201 wl_103 vdd gnd cell_6t
Xbit_r104_c201 bl_201 br_201 wl_104 vdd gnd cell_6t
Xbit_r105_c201 bl_201 br_201 wl_105 vdd gnd cell_6t
Xbit_r106_c201 bl_201 br_201 wl_106 vdd gnd cell_6t
Xbit_r107_c201 bl_201 br_201 wl_107 vdd gnd cell_6t
Xbit_r108_c201 bl_201 br_201 wl_108 vdd gnd cell_6t
Xbit_r109_c201 bl_201 br_201 wl_109 vdd gnd cell_6t
Xbit_r110_c201 bl_201 br_201 wl_110 vdd gnd cell_6t
Xbit_r111_c201 bl_201 br_201 wl_111 vdd gnd cell_6t
Xbit_r112_c201 bl_201 br_201 wl_112 vdd gnd cell_6t
Xbit_r113_c201 bl_201 br_201 wl_113 vdd gnd cell_6t
Xbit_r114_c201 bl_201 br_201 wl_114 vdd gnd cell_6t
Xbit_r115_c201 bl_201 br_201 wl_115 vdd gnd cell_6t
Xbit_r116_c201 bl_201 br_201 wl_116 vdd gnd cell_6t
Xbit_r117_c201 bl_201 br_201 wl_117 vdd gnd cell_6t
Xbit_r118_c201 bl_201 br_201 wl_118 vdd gnd cell_6t
Xbit_r119_c201 bl_201 br_201 wl_119 vdd gnd cell_6t
Xbit_r120_c201 bl_201 br_201 wl_120 vdd gnd cell_6t
Xbit_r121_c201 bl_201 br_201 wl_121 vdd gnd cell_6t
Xbit_r122_c201 bl_201 br_201 wl_122 vdd gnd cell_6t
Xbit_r123_c201 bl_201 br_201 wl_123 vdd gnd cell_6t
Xbit_r124_c201 bl_201 br_201 wl_124 vdd gnd cell_6t
Xbit_r125_c201 bl_201 br_201 wl_125 vdd gnd cell_6t
Xbit_r126_c201 bl_201 br_201 wl_126 vdd gnd cell_6t
Xbit_r127_c201 bl_201 br_201 wl_127 vdd gnd cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd cell_6t
Xbit_r1_c202 bl_202 br_202 wl_1 vdd gnd cell_6t
Xbit_r2_c202 bl_202 br_202 wl_2 vdd gnd cell_6t
Xbit_r3_c202 bl_202 br_202 wl_3 vdd gnd cell_6t
Xbit_r4_c202 bl_202 br_202 wl_4 vdd gnd cell_6t
Xbit_r5_c202 bl_202 br_202 wl_5 vdd gnd cell_6t
Xbit_r6_c202 bl_202 br_202 wl_6 vdd gnd cell_6t
Xbit_r7_c202 bl_202 br_202 wl_7 vdd gnd cell_6t
Xbit_r8_c202 bl_202 br_202 wl_8 vdd gnd cell_6t
Xbit_r9_c202 bl_202 br_202 wl_9 vdd gnd cell_6t
Xbit_r10_c202 bl_202 br_202 wl_10 vdd gnd cell_6t
Xbit_r11_c202 bl_202 br_202 wl_11 vdd gnd cell_6t
Xbit_r12_c202 bl_202 br_202 wl_12 vdd gnd cell_6t
Xbit_r13_c202 bl_202 br_202 wl_13 vdd gnd cell_6t
Xbit_r14_c202 bl_202 br_202 wl_14 vdd gnd cell_6t
Xbit_r15_c202 bl_202 br_202 wl_15 vdd gnd cell_6t
Xbit_r16_c202 bl_202 br_202 wl_16 vdd gnd cell_6t
Xbit_r17_c202 bl_202 br_202 wl_17 vdd gnd cell_6t
Xbit_r18_c202 bl_202 br_202 wl_18 vdd gnd cell_6t
Xbit_r19_c202 bl_202 br_202 wl_19 vdd gnd cell_6t
Xbit_r20_c202 bl_202 br_202 wl_20 vdd gnd cell_6t
Xbit_r21_c202 bl_202 br_202 wl_21 vdd gnd cell_6t
Xbit_r22_c202 bl_202 br_202 wl_22 vdd gnd cell_6t
Xbit_r23_c202 bl_202 br_202 wl_23 vdd gnd cell_6t
Xbit_r24_c202 bl_202 br_202 wl_24 vdd gnd cell_6t
Xbit_r25_c202 bl_202 br_202 wl_25 vdd gnd cell_6t
Xbit_r26_c202 bl_202 br_202 wl_26 vdd gnd cell_6t
Xbit_r27_c202 bl_202 br_202 wl_27 vdd gnd cell_6t
Xbit_r28_c202 bl_202 br_202 wl_28 vdd gnd cell_6t
Xbit_r29_c202 bl_202 br_202 wl_29 vdd gnd cell_6t
Xbit_r30_c202 bl_202 br_202 wl_30 vdd gnd cell_6t
Xbit_r31_c202 bl_202 br_202 wl_31 vdd gnd cell_6t
Xbit_r32_c202 bl_202 br_202 wl_32 vdd gnd cell_6t
Xbit_r33_c202 bl_202 br_202 wl_33 vdd gnd cell_6t
Xbit_r34_c202 bl_202 br_202 wl_34 vdd gnd cell_6t
Xbit_r35_c202 bl_202 br_202 wl_35 vdd gnd cell_6t
Xbit_r36_c202 bl_202 br_202 wl_36 vdd gnd cell_6t
Xbit_r37_c202 bl_202 br_202 wl_37 vdd gnd cell_6t
Xbit_r38_c202 bl_202 br_202 wl_38 vdd gnd cell_6t
Xbit_r39_c202 bl_202 br_202 wl_39 vdd gnd cell_6t
Xbit_r40_c202 bl_202 br_202 wl_40 vdd gnd cell_6t
Xbit_r41_c202 bl_202 br_202 wl_41 vdd gnd cell_6t
Xbit_r42_c202 bl_202 br_202 wl_42 vdd gnd cell_6t
Xbit_r43_c202 bl_202 br_202 wl_43 vdd gnd cell_6t
Xbit_r44_c202 bl_202 br_202 wl_44 vdd gnd cell_6t
Xbit_r45_c202 bl_202 br_202 wl_45 vdd gnd cell_6t
Xbit_r46_c202 bl_202 br_202 wl_46 vdd gnd cell_6t
Xbit_r47_c202 bl_202 br_202 wl_47 vdd gnd cell_6t
Xbit_r48_c202 bl_202 br_202 wl_48 vdd gnd cell_6t
Xbit_r49_c202 bl_202 br_202 wl_49 vdd gnd cell_6t
Xbit_r50_c202 bl_202 br_202 wl_50 vdd gnd cell_6t
Xbit_r51_c202 bl_202 br_202 wl_51 vdd gnd cell_6t
Xbit_r52_c202 bl_202 br_202 wl_52 vdd gnd cell_6t
Xbit_r53_c202 bl_202 br_202 wl_53 vdd gnd cell_6t
Xbit_r54_c202 bl_202 br_202 wl_54 vdd gnd cell_6t
Xbit_r55_c202 bl_202 br_202 wl_55 vdd gnd cell_6t
Xbit_r56_c202 bl_202 br_202 wl_56 vdd gnd cell_6t
Xbit_r57_c202 bl_202 br_202 wl_57 vdd gnd cell_6t
Xbit_r58_c202 bl_202 br_202 wl_58 vdd gnd cell_6t
Xbit_r59_c202 bl_202 br_202 wl_59 vdd gnd cell_6t
Xbit_r60_c202 bl_202 br_202 wl_60 vdd gnd cell_6t
Xbit_r61_c202 bl_202 br_202 wl_61 vdd gnd cell_6t
Xbit_r62_c202 bl_202 br_202 wl_62 vdd gnd cell_6t
Xbit_r63_c202 bl_202 br_202 wl_63 vdd gnd cell_6t
Xbit_r64_c202 bl_202 br_202 wl_64 vdd gnd cell_6t
Xbit_r65_c202 bl_202 br_202 wl_65 vdd gnd cell_6t
Xbit_r66_c202 bl_202 br_202 wl_66 vdd gnd cell_6t
Xbit_r67_c202 bl_202 br_202 wl_67 vdd gnd cell_6t
Xbit_r68_c202 bl_202 br_202 wl_68 vdd gnd cell_6t
Xbit_r69_c202 bl_202 br_202 wl_69 vdd gnd cell_6t
Xbit_r70_c202 bl_202 br_202 wl_70 vdd gnd cell_6t
Xbit_r71_c202 bl_202 br_202 wl_71 vdd gnd cell_6t
Xbit_r72_c202 bl_202 br_202 wl_72 vdd gnd cell_6t
Xbit_r73_c202 bl_202 br_202 wl_73 vdd gnd cell_6t
Xbit_r74_c202 bl_202 br_202 wl_74 vdd gnd cell_6t
Xbit_r75_c202 bl_202 br_202 wl_75 vdd gnd cell_6t
Xbit_r76_c202 bl_202 br_202 wl_76 vdd gnd cell_6t
Xbit_r77_c202 bl_202 br_202 wl_77 vdd gnd cell_6t
Xbit_r78_c202 bl_202 br_202 wl_78 vdd gnd cell_6t
Xbit_r79_c202 bl_202 br_202 wl_79 vdd gnd cell_6t
Xbit_r80_c202 bl_202 br_202 wl_80 vdd gnd cell_6t
Xbit_r81_c202 bl_202 br_202 wl_81 vdd gnd cell_6t
Xbit_r82_c202 bl_202 br_202 wl_82 vdd gnd cell_6t
Xbit_r83_c202 bl_202 br_202 wl_83 vdd gnd cell_6t
Xbit_r84_c202 bl_202 br_202 wl_84 vdd gnd cell_6t
Xbit_r85_c202 bl_202 br_202 wl_85 vdd gnd cell_6t
Xbit_r86_c202 bl_202 br_202 wl_86 vdd gnd cell_6t
Xbit_r87_c202 bl_202 br_202 wl_87 vdd gnd cell_6t
Xbit_r88_c202 bl_202 br_202 wl_88 vdd gnd cell_6t
Xbit_r89_c202 bl_202 br_202 wl_89 vdd gnd cell_6t
Xbit_r90_c202 bl_202 br_202 wl_90 vdd gnd cell_6t
Xbit_r91_c202 bl_202 br_202 wl_91 vdd gnd cell_6t
Xbit_r92_c202 bl_202 br_202 wl_92 vdd gnd cell_6t
Xbit_r93_c202 bl_202 br_202 wl_93 vdd gnd cell_6t
Xbit_r94_c202 bl_202 br_202 wl_94 vdd gnd cell_6t
Xbit_r95_c202 bl_202 br_202 wl_95 vdd gnd cell_6t
Xbit_r96_c202 bl_202 br_202 wl_96 vdd gnd cell_6t
Xbit_r97_c202 bl_202 br_202 wl_97 vdd gnd cell_6t
Xbit_r98_c202 bl_202 br_202 wl_98 vdd gnd cell_6t
Xbit_r99_c202 bl_202 br_202 wl_99 vdd gnd cell_6t
Xbit_r100_c202 bl_202 br_202 wl_100 vdd gnd cell_6t
Xbit_r101_c202 bl_202 br_202 wl_101 vdd gnd cell_6t
Xbit_r102_c202 bl_202 br_202 wl_102 vdd gnd cell_6t
Xbit_r103_c202 bl_202 br_202 wl_103 vdd gnd cell_6t
Xbit_r104_c202 bl_202 br_202 wl_104 vdd gnd cell_6t
Xbit_r105_c202 bl_202 br_202 wl_105 vdd gnd cell_6t
Xbit_r106_c202 bl_202 br_202 wl_106 vdd gnd cell_6t
Xbit_r107_c202 bl_202 br_202 wl_107 vdd gnd cell_6t
Xbit_r108_c202 bl_202 br_202 wl_108 vdd gnd cell_6t
Xbit_r109_c202 bl_202 br_202 wl_109 vdd gnd cell_6t
Xbit_r110_c202 bl_202 br_202 wl_110 vdd gnd cell_6t
Xbit_r111_c202 bl_202 br_202 wl_111 vdd gnd cell_6t
Xbit_r112_c202 bl_202 br_202 wl_112 vdd gnd cell_6t
Xbit_r113_c202 bl_202 br_202 wl_113 vdd gnd cell_6t
Xbit_r114_c202 bl_202 br_202 wl_114 vdd gnd cell_6t
Xbit_r115_c202 bl_202 br_202 wl_115 vdd gnd cell_6t
Xbit_r116_c202 bl_202 br_202 wl_116 vdd gnd cell_6t
Xbit_r117_c202 bl_202 br_202 wl_117 vdd gnd cell_6t
Xbit_r118_c202 bl_202 br_202 wl_118 vdd gnd cell_6t
Xbit_r119_c202 bl_202 br_202 wl_119 vdd gnd cell_6t
Xbit_r120_c202 bl_202 br_202 wl_120 vdd gnd cell_6t
Xbit_r121_c202 bl_202 br_202 wl_121 vdd gnd cell_6t
Xbit_r122_c202 bl_202 br_202 wl_122 vdd gnd cell_6t
Xbit_r123_c202 bl_202 br_202 wl_123 vdd gnd cell_6t
Xbit_r124_c202 bl_202 br_202 wl_124 vdd gnd cell_6t
Xbit_r125_c202 bl_202 br_202 wl_125 vdd gnd cell_6t
Xbit_r126_c202 bl_202 br_202 wl_126 vdd gnd cell_6t
Xbit_r127_c202 bl_202 br_202 wl_127 vdd gnd cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd cell_6t
Xbit_r1_c203 bl_203 br_203 wl_1 vdd gnd cell_6t
Xbit_r2_c203 bl_203 br_203 wl_2 vdd gnd cell_6t
Xbit_r3_c203 bl_203 br_203 wl_3 vdd gnd cell_6t
Xbit_r4_c203 bl_203 br_203 wl_4 vdd gnd cell_6t
Xbit_r5_c203 bl_203 br_203 wl_5 vdd gnd cell_6t
Xbit_r6_c203 bl_203 br_203 wl_6 vdd gnd cell_6t
Xbit_r7_c203 bl_203 br_203 wl_7 vdd gnd cell_6t
Xbit_r8_c203 bl_203 br_203 wl_8 vdd gnd cell_6t
Xbit_r9_c203 bl_203 br_203 wl_9 vdd gnd cell_6t
Xbit_r10_c203 bl_203 br_203 wl_10 vdd gnd cell_6t
Xbit_r11_c203 bl_203 br_203 wl_11 vdd gnd cell_6t
Xbit_r12_c203 bl_203 br_203 wl_12 vdd gnd cell_6t
Xbit_r13_c203 bl_203 br_203 wl_13 vdd gnd cell_6t
Xbit_r14_c203 bl_203 br_203 wl_14 vdd gnd cell_6t
Xbit_r15_c203 bl_203 br_203 wl_15 vdd gnd cell_6t
Xbit_r16_c203 bl_203 br_203 wl_16 vdd gnd cell_6t
Xbit_r17_c203 bl_203 br_203 wl_17 vdd gnd cell_6t
Xbit_r18_c203 bl_203 br_203 wl_18 vdd gnd cell_6t
Xbit_r19_c203 bl_203 br_203 wl_19 vdd gnd cell_6t
Xbit_r20_c203 bl_203 br_203 wl_20 vdd gnd cell_6t
Xbit_r21_c203 bl_203 br_203 wl_21 vdd gnd cell_6t
Xbit_r22_c203 bl_203 br_203 wl_22 vdd gnd cell_6t
Xbit_r23_c203 bl_203 br_203 wl_23 vdd gnd cell_6t
Xbit_r24_c203 bl_203 br_203 wl_24 vdd gnd cell_6t
Xbit_r25_c203 bl_203 br_203 wl_25 vdd gnd cell_6t
Xbit_r26_c203 bl_203 br_203 wl_26 vdd gnd cell_6t
Xbit_r27_c203 bl_203 br_203 wl_27 vdd gnd cell_6t
Xbit_r28_c203 bl_203 br_203 wl_28 vdd gnd cell_6t
Xbit_r29_c203 bl_203 br_203 wl_29 vdd gnd cell_6t
Xbit_r30_c203 bl_203 br_203 wl_30 vdd gnd cell_6t
Xbit_r31_c203 bl_203 br_203 wl_31 vdd gnd cell_6t
Xbit_r32_c203 bl_203 br_203 wl_32 vdd gnd cell_6t
Xbit_r33_c203 bl_203 br_203 wl_33 vdd gnd cell_6t
Xbit_r34_c203 bl_203 br_203 wl_34 vdd gnd cell_6t
Xbit_r35_c203 bl_203 br_203 wl_35 vdd gnd cell_6t
Xbit_r36_c203 bl_203 br_203 wl_36 vdd gnd cell_6t
Xbit_r37_c203 bl_203 br_203 wl_37 vdd gnd cell_6t
Xbit_r38_c203 bl_203 br_203 wl_38 vdd gnd cell_6t
Xbit_r39_c203 bl_203 br_203 wl_39 vdd gnd cell_6t
Xbit_r40_c203 bl_203 br_203 wl_40 vdd gnd cell_6t
Xbit_r41_c203 bl_203 br_203 wl_41 vdd gnd cell_6t
Xbit_r42_c203 bl_203 br_203 wl_42 vdd gnd cell_6t
Xbit_r43_c203 bl_203 br_203 wl_43 vdd gnd cell_6t
Xbit_r44_c203 bl_203 br_203 wl_44 vdd gnd cell_6t
Xbit_r45_c203 bl_203 br_203 wl_45 vdd gnd cell_6t
Xbit_r46_c203 bl_203 br_203 wl_46 vdd gnd cell_6t
Xbit_r47_c203 bl_203 br_203 wl_47 vdd gnd cell_6t
Xbit_r48_c203 bl_203 br_203 wl_48 vdd gnd cell_6t
Xbit_r49_c203 bl_203 br_203 wl_49 vdd gnd cell_6t
Xbit_r50_c203 bl_203 br_203 wl_50 vdd gnd cell_6t
Xbit_r51_c203 bl_203 br_203 wl_51 vdd gnd cell_6t
Xbit_r52_c203 bl_203 br_203 wl_52 vdd gnd cell_6t
Xbit_r53_c203 bl_203 br_203 wl_53 vdd gnd cell_6t
Xbit_r54_c203 bl_203 br_203 wl_54 vdd gnd cell_6t
Xbit_r55_c203 bl_203 br_203 wl_55 vdd gnd cell_6t
Xbit_r56_c203 bl_203 br_203 wl_56 vdd gnd cell_6t
Xbit_r57_c203 bl_203 br_203 wl_57 vdd gnd cell_6t
Xbit_r58_c203 bl_203 br_203 wl_58 vdd gnd cell_6t
Xbit_r59_c203 bl_203 br_203 wl_59 vdd gnd cell_6t
Xbit_r60_c203 bl_203 br_203 wl_60 vdd gnd cell_6t
Xbit_r61_c203 bl_203 br_203 wl_61 vdd gnd cell_6t
Xbit_r62_c203 bl_203 br_203 wl_62 vdd gnd cell_6t
Xbit_r63_c203 bl_203 br_203 wl_63 vdd gnd cell_6t
Xbit_r64_c203 bl_203 br_203 wl_64 vdd gnd cell_6t
Xbit_r65_c203 bl_203 br_203 wl_65 vdd gnd cell_6t
Xbit_r66_c203 bl_203 br_203 wl_66 vdd gnd cell_6t
Xbit_r67_c203 bl_203 br_203 wl_67 vdd gnd cell_6t
Xbit_r68_c203 bl_203 br_203 wl_68 vdd gnd cell_6t
Xbit_r69_c203 bl_203 br_203 wl_69 vdd gnd cell_6t
Xbit_r70_c203 bl_203 br_203 wl_70 vdd gnd cell_6t
Xbit_r71_c203 bl_203 br_203 wl_71 vdd gnd cell_6t
Xbit_r72_c203 bl_203 br_203 wl_72 vdd gnd cell_6t
Xbit_r73_c203 bl_203 br_203 wl_73 vdd gnd cell_6t
Xbit_r74_c203 bl_203 br_203 wl_74 vdd gnd cell_6t
Xbit_r75_c203 bl_203 br_203 wl_75 vdd gnd cell_6t
Xbit_r76_c203 bl_203 br_203 wl_76 vdd gnd cell_6t
Xbit_r77_c203 bl_203 br_203 wl_77 vdd gnd cell_6t
Xbit_r78_c203 bl_203 br_203 wl_78 vdd gnd cell_6t
Xbit_r79_c203 bl_203 br_203 wl_79 vdd gnd cell_6t
Xbit_r80_c203 bl_203 br_203 wl_80 vdd gnd cell_6t
Xbit_r81_c203 bl_203 br_203 wl_81 vdd gnd cell_6t
Xbit_r82_c203 bl_203 br_203 wl_82 vdd gnd cell_6t
Xbit_r83_c203 bl_203 br_203 wl_83 vdd gnd cell_6t
Xbit_r84_c203 bl_203 br_203 wl_84 vdd gnd cell_6t
Xbit_r85_c203 bl_203 br_203 wl_85 vdd gnd cell_6t
Xbit_r86_c203 bl_203 br_203 wl_86 vdd gnd cell_6t
Xbit_r87_c203 bl_203 br_203 wl_87 vdd gnd cell_6t
Xbit_r88_c203 bl_203 br_203 wl_88 vdd gnd cell_6t
Xbit_r89_c203 bl_203 br_203 wl_89 vdd gnd cell_6t
Xbit_r90_c203 bl_203 br_203 wl_90 vdd gnd cell_6t
Xbit_r91_c203 bl_203 br_203 wl_91 vdd gnd cell_6t
Xbit_r92_c203 bl_203 br_203 wl_92 vdd gnd cell_6t
Xbit_r93_c203 bl_203 br_203 wl_93 vdd gnd cell_6t
Xbit_r94_c203 bl_203 br_203 wl_94 vdd gnd cell_6t
Xbit_r95_c203 bl_203 br_203 wl_95 vdd gnd cell_6t
Xbit_r96_c203 bl_203 br_203 wl_96 vdd gnd cell_6t
Xbit_r97_c203 bl_203 br_203 wl_97 vdd gnd cell_6t
Xbit_r98_c203 bl_203 br_203 wl_98 vdd gnd cell_6t
Xbit_r99_c203 bl_203 br_203 wl_99 vdd gnd cell_6t
Xbit_r100_c203 bl_203 br_203 wl_100 vdd gnd cell_6t
Xbit_r101_c203 bl_203 br_203 wl_101 vdd gnd cell_6t
Xbit_r102_c203 bl_203 br_203 wl_102 vdd gnd cell_6t
Xbit_r103_c203 bl_203 br_203 wl_103 vdd gnd cell_6t
Xbit_r104_c203 bl_203 br_203 wl_104 vdd gnd cell_6t
Xbit_r105_c203 bl_203 br_203 wl_105 vdd gnd cell_6t
Xbit_r106_c203 bl_203 br_203 wl_106 vdd gnd cell_6t
Xbit_r107_c203 bl_203 br_203 wl_107 vdd gnd cell_6t
Xbit_r108_c203 bl_203 br_203 wl_108 vdd gnd cell_6t
Xbit_r109_c203 bl_203 br_203 wl_109 vdd gnd cell_6t
Xbit_r110_c203 bl_203 br_203 wl_110 vdd gnd cell_6t
Xbit_r111_c203 bl_203 br_203 wl_111 vdd gnd cell_6t
Xbit_r112_c203 bl_203 br_203 wl_112 vdd gnd cell_6t
Xbit_r113_c203 bl_203 br_203 wl_113 vdd gnd cell_6t
Xbit_r114_c203 bl_203 br_203 wl_114 vdd gnd cell_6t
Xbit_r115_c203 bl_203 br_203 wl_115 vdd gnd cell_6t
Xbit_r116_c203 bl_203 br_203 wl_116 vdd gnd cell_6t
Xbit_r117_c203 bl_203 br_203 wl_117 vdd gnd cell_6t
Xbit_r118_c203 bl_203 br_203 wl_118 vdd gnd cell_6t
Xbit_r119_c203 bl_203 br_203 wl_119 vdd gnd cell_6t
Xbit_r120_c203 bl_203 br_203 wl_120 vdd gnd cell_6t
Xbit_r121_c203 bl_203 br_203 wl_121 vdd gnd cell_6t
Xbit_r122_c203 bl_203 br_203 wl_122 vdd gnd cell_6t
Xbit_r123_c203 bl_203 br_203 wl_123 vdd gnd cell_6t
Xbit_r124_c203 bl_203 br_203 wl_124 vdd gnd cell_6t
Xbit_r125_c203 bl_203 br_203 wl_125 vdd gnd cell_6t
Xbit_r126_c203 bl_203 br_203 wl_126 vdd gnd cell_6t
Xbit_r127_c203 bl_203 br_203 wl_127 vdd gnd cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd cell_6t
Xbit_r1_c204 bl_204 br_204 wl_1 vdd gnd cell_6t
Xbit_r2_c204 bl_204 br_204 wl_2 vdd gnd cell_6t
Xbit_r3_c204 bl_204 br_204 wl_3 vdd gnd cell_6t
Xbit_r4_c204 bl_204 br_204 wl_4 vdd gnd cell_6t
Xbit_r5_c204 bl_204 br_204 wl_5 vdd gnd cell_6t
Xbit_r6_c204 bl_204 br_204 wl_6 vdd gnd cell_6t
Xbit_r7_c204 bl_204 br_204 wl_7 vdd gnd cell_6t
Xbit_r8_c204 bl_204 br_204 wl_8 vdd gnd cell_6t
Xbit_r9_c204 bl_204 br_204 wl_9 vdd gnd cell_6t
Xbit_r10_c204 bl_204 br_204 wl_10 vdd gnd cell_6t
Xbit_r11_c204 bl_204 br_204 wl_11 vdd gnd cell_6t
Xbit_r12_c204 bl_204 br_204 wl_12 vdd gnd cell_6t
Xbit_r13_c204 bl_204 br_204 wl_13 vdd gnd cell_6t
Xbit_r14_c204 bl_204 br_204 wl_14 vdd gnd cell_6t
Xbit_r15_c204 bl_204 br_204 wl_15 vdd gnd cell_6t
Xbit_r16_c204 bl_204 br_204 wl_16 vdd gnd cell_6t
Xbit_r17_c204 bl_204 br_204 wl_17 vdd gnd cell_6t
Xbit_r18_c204 bl_204 br_204 wl_18 vdd gnd cell_6t
Xbit_r19_c204 bl_204 br_204 wl_19 vdd gnd cell_6t
Xbit_r20_c204 bl_204 br_204 wl_20 vdd gnd cell_6t
Xbit_r21_c204 bl_204 br_204 wl_21 vdd gnd cell_6t
Xbit_r22_c204 bl_204 br_204 wl_22 vdd gnd cell_6t
Xbit_r23_c204 bl_204 br_204 wl_23 vdd gnd cell_6t
Xbit_r24_c204 bl_204 br_204 wl_24 vdd gnd cell_6t
Xbit_r25_c204 bl_204 br_204 wl_25 vdd gnd cell_6t
Xbit_r26_c204 bl_204 br_204 wl_26 vdd gnd cell_6t
Xbit_r27_c204 bl_204 br_204 wl_27 vdd gnd cell_6t
Xbit_r28_c204 bl_204 br_204 wl_28 vdd gnd cell_6t
Xbit_r29_c204 bl_204 br_204 wl_29 vdd gnd cell_6t
Xbit_r30_c204 bl_204 br_204 wl_30 vdd gnd cell_6t
Xbit_r31_c204 bl_204 br_204 wl_31 vdd gnd cell_6t
Xbit_r32_c204 bl_204 br_204 wl_32 vdd gnd cell_6t
Xbit_r33_c204 bl_204 br_204 wl_33 vdd gnd cell_6t
Xbit_r34_c204 bl_204 br_204 wl_34 vdd gnd cell_6t
Xbit_r35_c204 bl_204 br_204 wl_35 vdd gnd cell_6t
Xbit_r36_c204 bl_204 br_204 wl_36 vdd gnd cell_6t
Xbit_r37_c204 bl_204 br_204 wl_37 vdd gnd cell_6t
Xbit_r38_c204 bl_204 br_204 wl_38 vdd gnd cell_6t
Xbit_r39_c204 bl_204 br_204 wl_39 vdd gnd cell_6t
Xbit_r40_c204 bl_204 br_204 wl_40 vdd gnd cell_6t
Xbit_r41_c204 bl_204 br_204 wl_41 vdd gnd cell_6t
Xbit_r42_c204 bl_204 br_204 wl_42 vdd gnd cell_6t
Xbit_r43_c204 bl_204 br_204 wl_43 vdd gnd cell_6t
Xbit_r44_c204 bl_204 br_204 wl_44 vdd gnd cell_6t
Xbit_r45_c204 bl_204 br_204 wl_45 vdd gnd cell_6t
Xbit_r46_c204 bl_204 br_204 wl_46 vdd gnd cell_6t
Xbit_r47_c204 bl_204 br_204 wl_47 vdd gnd cell_6t
Xbit_r48_c204 bl_204 br_204 wl_48 vdd gnd cell_6t
Xbit_r49_c204 bl_204 br_204 wl_49 vdd gnd cell_6t
Xbit_r50_c204 bl_204 br_204 wl_50 vdd gnd cell_6t
Xbit_r51_c204 bl_204 br_204 wl_51 vdd gnd cell_6t
Xbit_r52_c204 bl_204 br_204 wl_52 vdd gnd cell_6t
Xbit_r53_c204 bl_204 br_204 wl_53 vdd gnd cell_6t
Xbit_r54_c204 bl_204 br_204 wl_54 vdd gnd cell_6t
Xbit_r55_c204 bl_204 br_204 wl_55 vdd gnd cell_6t
Xbit_r56_c204 bl_204 br_204 wl_56 vdd gnd cell_6t
Xbit_r57_c204 bl_204 br_204 wl_57 vdd gnd cell_6t
Xbit_r58_c204 bl_204 br_204 wl_58 vdd gnd cell_6t
Xbit_r59_c204 bl_204 br_204 wl_59 vdd gnd cell_6t
Xbit_r60_c204 bl_204 br_204 wl_60 vdd gnd cell_6t
Xbit_r61_c204 bl_204 br_204 wl_61 vdd gnd cell_6t
Xbit_r62_c204 bl_204 br_204 wl_62 vdd gnd cell_6t
Xbit_r63_c204 bl_204 br_204 wl_63 vdd gnd cell_6t
Xbit_r64_c204 bl_204 br_204 wl_64 vdd gnd cell_6t
Xbit_r65_c204 bl_204 br_204 wl_65 vdd gnd cell_6t
Xbit_r66_c204 bl_204 br_204 wl_66 vdd gnd cell_6t
Xbit_r67_c204 bl_204 br_204 wl_67 vdd gnd cell_6t
Xbit_r68_c204 bl_204 br_204 wl_68 vdd gnd cell_6t
Xbit_r69_c204 bl_204 br_204 wl_69 vdd gnd cell_6t
Xbit_r70_c204 bl_204 br_204 wl_70 vdd gnd cell_6t
Xbit_r71_c204 bl_204 br_204 wl_71 vdd gnd cell_6t
Xbit_r72_c204 bl_204 br_204 wl_72 vdd gnd cell_6t
Xbit_r73_c204 bl_204 br_204 wl_73 vdd gnd cell_6t
Xbit_r74_c204 bl_204 br_204 wl_74 vdd gnd cell_6t
Xbit_r75_c204 bl_204 br_204 wl_75 vdd gnd cell_6t
Xbit_r76_c204 bl_204 br_204 wl_76 vdd gnd cell_6t
Xbit_r77_c204 bl_204 br_204 wl_77 vdd gnd cell_6t
Xbit_r78_c204 bl_204 br_204 wl_78 vdd gnd cell_6t
Xbit_r79_c204 bl_204 br_204 wl_79 vdd gnd cell_6t
Xbit_r80_c204 bl_204 br_204 wl_80 vdd gnd cell_6t
Xbit_r81_c204 bl_204 br_204 wl_81 vdd gnd cell_6t
Xbit_r82_c204 bl_204 br_204 wl_82 vdd gnd cell_6t
Xbit_r83_c204 bl_204 br_204 wl_83 vdd gnd cell_6t
Xbit_r84_c204 bl_204 br_204 wl_84 vdd gnd cell_6t
Xbit_r85_c204 bl_204 br_204 wl_85 vdd gnd cell_6t
Xbit_r86_c204 bl_204 br_204 wl_86 vdd gnd cell_6t
Xbit_r87_c204 bl_204 br_204 wl_87 vdd gnd cell_6t
Xbit_r88_c204 bl_204 br_204 wl_88 vdd gnd cell_6t
Xbit_r89_c204 bl_204 br_204 wl_89 vdd gnd cell_6t
Xbit_r90_c204 bl_204 br_204 wl_90 vdd gnd cell_6t
Xbit_r91_c204 bl_204 br_204 wl_91 vdd gnd cell_6t
Xbit_r92_c204 bl_204 br_204 wl_92 vdd gnd cell_6t
Xbit_r93_c204 bl_204 br_204 wl_93 vdd gnd cell_6t
Xbit_r94_c204 bl_204 br_204 wl_94 vdd gnd cell_6t
Xbit_r95_c204 bl_204 br_204 wl_95 vdd gnd cell_6t
Xbit_r96_c204 bl_204 br_204 wl_96 vdd gnd cell_6t
Xbit_r97_c204 bl_204 br_204 wl_97 vdd gnd cell_6t
Xbit_r98_c204 bl_204 br_204 wl_98 vdd gnd cell_6t
Xbit_r99_c204 bl_204 br_204 wl_99 vdd gnd cell_6t
Xbit_r100_c204 bl_204 br_204 wl_100 vdd gnd cell_6t
Xbit_r101_c204 bl_204 br_204 wl_101 vdd gnd cell_6t
Xbit_r102_c204 bl_204 br_204 wl_102 vdd gnd cell_6t
Xbit_r103_c204 bl_204 br_204 wl_103 vdd gnd cell_6t
Xbit_r104_c204 bl_204 br_204 wl_104 vdd gnd cell_6t
Xbit_r105_c204 bl_204 br_204 wl_105 vdd gnd cell_6t
Xbit_r106_c204 bl_204 br_204 wl_106 vdd gnd cell_6t
Xbit_r107_c204 bl_204 br_204 wl_107 vdd gnd cell_6t
Xbit_r108_c204 bl_204 br_204 wl_108 vdd gnd cell_6t
Xbit_r109_c204 bl_204 br_204 wl_109 vdd gnd cell_6t
Xbit_r110_c204 bl_204 br_204 wl_110 vdd gnd cell_6t
Xbit_r111_c204 bl_204 br_204 wl_111 vdd gnd cell_6t
Xbit_r112_c204 bl_204 br_204 wl_112 vdd gnd cell_6t
Xbit_r113_c204 bl_204 br_204 wl_113 vdd gnd cell_6t
Xbit_r114_c204 bl_204 br_204 wl_114 vdd gnd cell_6t
Xbit_r115_c204 bl_204 br_204 wl_115 vdd gnd cell_6t
Xbit_r116_c204 bl_204 br_204 wl_116 vdd gnd cell_6t
Xbit_r117_c204 bl_204 br_204 wl_117 vdd gnd cell_6t
Xbit_r118_c204 bl_204 br_204 wl_118 vdd gnd cell_6t
Xbit_r119_c204 bl_204 br_204 wl_119 vdd gnd cell_6t
Xbit_r120_c204 bl_204 br_204 wl_120 vdd gnd cell_6t
Xbit_r121_c204 bl_204 br_204 wl_121 vdd gnd cell_6t
Xbit_r122_c204 bl_204 br_204 wl_122 vdd gnd cell_6t
Xbit_r123_c204 bl_204 br_204 wl_123 vdd gnd cell_6t
Xbit_r124_c204 bl_204 br_204 wl_124 vdd gnd cell_6t
Xbit_r125_c204 bl_204 br_204 wl_125 vdd gnd cell_6t
Xbit_r126_c204 bl_204 br_204 wl_126 vdd gnd cell_6t
Xbit_r127_c204 bl_204 br_204 wl_127 vdd gnd cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd cell_6t
Xbit_r1_c205 bl_205 br_205 wl_1 vdd gnd cell_6t
Xbit_r2_c205 bl_205 br_205 wl_2 vdd gnd cell_6t
Xbit_r3_c205 bl_205 br_205 wl_3 vdd gnd cell_6t
Xbit_r4_c205 bl_205 br_205 wl_4 vdd gnd cell_6t
Xbit_r5_c205 bl_205 br_205 wl_5 vdd gnd cell_6t
Xbit_r6_c205 bl_205 br_205 wl_6 vdd gnd cell_6t
Xbit_r7_c205 bl_205 br_205 wl_7 vdd gnd cell_6t
Xbit_r8_c205 bl_205 br_205 wl_8 vdd gnd cell_6t
Xbit_r9_c205 bl_205 br_205 wl_9 vdd gnd cell_6t
Xbit_r10_c205 bl_205 br_205 wl_10 vdd gnd cell_6t
Xbit_r11_c205 bl_205 br_205 wl_11 vdd gnd cell_6t
Xbit_r12_c205 bl_205 br_205 wl_12 vdd gnd cell_6t
Xbit_r13_c205 bl_205 br_205 wl_13 vdd gnd cell_6t
Xbit_r14_c205 bl_205 br_205 wl_14 vdd gnd cell_6t
Xbit_r15_c205 bl_205 br_205 wl_15 vdd gnd cell_6t
Xbit_r16_c205 bl_205 br_205 wl_16 vdd gnd cell_6t
Xbit_r17_c205 bl_205 br_205 wl_17 vdd gnd cell_6t
Xbit_r18_c205 bl_205 br_205 wl_18 vdd gnd cell_6t
Xbit_r19_c205 bl_205 br_205 wl_19 vdd gnd cell_6t
Xbit_r20_c205 bl_205 br_205 wl_20 vdd gnd cell_6t
Xbit_r21_c205 bl_205 br_205 wl_21 vdd gnd cell_6t
Xbit_r22_c205 bl_205 br_205 wl_22 vdd gnd cell_6t
Xbit_r23_c205 bl_205 br_205 wl_23 vdd gnd cell_6t
Xbit_r24_c205 bl_205 br_205 wl_24 vdd gnd cell_6t
Xbit_r25_c205 bl_205 br_205 wl_25 vdd gnd cell_6t
Xbit_r26_c205 bl_205 br_205 wl_26 vdd gnd cell_6t
Xbit_r27_c205 bl_205 br_205 wl_27 vdd gnd cell_6t
Xbit_r28_c205 bl_205 br_205 wl_28 vdd gnd cell_6t
Xbit_r29_c205 bl_205 br_205 wl_29 vdd gnd cell_6t
Xbit_r30_c205 bl_205 br_205 wl_30 vdd gnd cell_6t
Xbit_r31_c205 bl_205 br_205 wl_31 vdd gnd cell_6t
Xbit_r32_c205 bl_205 br_205 wl_32 vdd gnd cell_6t
Xbit_r33_c205 bl_205 br_205 wl_33 vdd gnd cell_6t
Xbit_r34_c205 bl_205 br_205 wl_34 vdd gnd cell_6t
Xbit_r35_c205 bl_205 br_205 wl_35 vdd gnd cell_6t
Xbit_r36_c205 bl_205 br_205 wl_36 vdd gnd cell_6t
Xbit_r37_c205 bl_205 br_205 wl_37 vdd gnd cell_6t
Xbit_r38_c205 bl_205 br_205 wl_38 vdd gnd cell_6t
Xbit_r39_c205 bl_205 br_205 wl_39 vdd gnd cell_6t
Xbit_r40_c205 bl_205 br_205 wl_40 vdd gnd cell_6t
Xbit_r41_c205 bl_205 br_205 wl_41 vdd gnd cell_6t
Xbit_r42_c205 bl_205 br_205 wl_42 vdd gnd cell_6t
Xbit_r43_c205 bl_205 br_205 wl_43 vdd gnd cell_6t
Xbit_r44_c205 bl_205 br_205 wl_44 vdd gnd cell_6t
Xbit_r45_c205 bl_205 br_205 wl_45 vdd gnd cell_6t
Xbit_r46_c205 bl_205 br_205 wl_46 vdd gnd cell_6t
Xbit_r47_c205 bl_205 br_205 wl_47 vdd gnd cell_6t
Xbit_r48_c205 bl_205 br_205 wl_48 vdd gnd cell_6t
Xbit_r49_c205 bl_205 br_205 wl_49 vdd gnd cell_6t
Xbit_r50_c205 bl_205 br_205 wl_50 vdd gnd cell_6t
Xbit_r51_c205 bl_205 br_205 wl_51 vdd gnd cell_6t
Xbit_r52_c205 bl_205 br_205 wl_52 vdd gnd cell_6t
Xbit_r53_c205 bl_205 br_205 wl_53 vdd gnd cell_6t
Xbit_r54_c205 bl_205 br_205 wl_54 vdd gnd cell_6t
Xbit_r55_c205 bl_205 br_205 wl_55 vdd gnd cell_6t
Xbit_r56_c205 bl_205 br_205 wl_56 vdd gnd cell_6t
Xbit_r57_c205 bl_205 br_205 wl_57 vdd gnd cell_6t
Xbit_r58_c205 bl_205 br_205 wl_58 vdd gnd cell_6t
Xbit_r59_c205 bl_205 br_205 wl_59 vdd gnd cell_6t
Xbit_r60_c205 bl_205 br_205 wl_60 vdd gnd cell_6t
Xbit_r61_c205 bl_205 br_205 wl_61 vdd gnd cell_6t
Xbit_r62_c205 bl_205 br_205 wl_62 vdd gnd cell_6t
Xbit_r63_c205 bl_205 br_205 wl_63 vdd gnd cell_6t
Xbit_r64_c205 bl_205 br_205 wl_64 vdd gnd cell_6t
Xbit_r65_c205 bl_205 br_205 wl_65 vdd gnd cell_6t
Xbit_r66_c205 bl_205 br_205 wl_66 vdd gnd cell_6t
Xbit_r67_c205 bl_205 br_205 wl_67 vdd gnd cell_6t
Xbit_r68_c205 bl_205 br_205 wl_68 vdd gnd cell_6t
Xbit_r69_c205 bl_205 br_205 wl_69 vdd gnd cell_6t
Xbit_r70_c205 bl_205 br_205 wl_70 vdd gnd cell_6t
Xbit_r71_c205 bl_205 br_205 wl_71 vdd gnd cell_6t
Xbit_r72_c205 bl_205 br_205 wl_72 vdd gnd cell_6t
Xbit_r73_c205 bl_205 br_205 wl_73 vdd gnd cell_6t
Xbit_r74_c205 bl_205 br_205 wl_74 vdd gnd cell_6t
Xbit_r75_c205 bl_205 br_205 wl_75 vdd gnd cell_6t
Xbit_r76_c205 bl_205 br_205 wl_76 vdd gnd cell_6t
Xbit_r77_c205 bl_205 br_205 wl_77 vdd gnd cell_6t
Xbit_r78_c205 bl_205 br_205 wl_78 vdd gnd cell_6t
Xbit_r79_c205 bl_205 br_205 wl_79 vdd gnd cell_6t
Xbit_r80_c205 bl_205 br_205 wl_80 vdd gnd cell_6t
Xbit_r81_c205 bl_205 br_205 wl_81 vdd gnd cell_6t
Xbit_r82_c205 bl_205 br_205 wl_82 vdd gnd cell_6t
Xbit_r83_c205 bl_205 br_205 wl_83 vdd gnd cell_6t
Xbit_r84_c205 bl_205 br_205 wl_84 vdd gnd cell_6t
Xbit_r85_c205 bl_205 br_205 wl_85 vdd gnd cell_6t
Xbit_r86_c205 bl_205 br_205 wl_86 vdd gnd cell_6t
Xbit_r87_c205 bl_205 br_205 wl_87 vdd gnd cell_6t
Xbit_r88_c205 bl_205 br_205 wl_88 vdd gnd cell_6t
Xbit_r89_c205 bl_205 br_205 wl_89 vdd gnd cell_6t
Xbit_r90_c205 bl_205 br_205 wl_90 vdd gnd cell_6t
Xbit_r91_c205 bl_205 br_205 wl_91 vdd gnd cell_6t
Xbit_r92_c205 bl_205 br_205 wl_92 vdd gnd cell_6t
Xbit_r93_c205 bl_205 br_205 wl_93 vdd gnd cell_6t
Xbit_r94_c205 bl_205 br_205 wl_94 vdd gnd cell_6t
Xbit_r95_c205 bl_205 br_205 wl_95 vdd gnd cell_6t
Xbit_r96_c205 bl_205 br_205 wl_96 vdd gnd cell_6t
Xbit_r97_c205 bl_205 br_205 wl_97 vdd gnd cell_6t
Xbit_r98_c205 bl_205 br_205 wl_98 vdd gnd cell_6t
Xbit_r99_c205 bl_205 br_205 wl_99 vdd gnd cell_6t
Xbit_r100_c205 bl_205 br_205 wl_100 vdd gnd cell_6t
Xbit_r101_c205 bl_205 br_205 wl_101 vdd gnd cell_6t
Xbit_r102_c205 bl_205 br_205 wl_102 vdd gnd cell_6t
Xbit_r103_c205 bl_205 br_205 wl_103 vdd gnd cell_6t
Xbit_r104_c205 bl_205 br_205 wl_104 vdd gnd cell_6t
Xbit_r105_c205 bl_205 br_205 wl_105 vdd gnd cell_6t
Xbit_r106_c205 bl_205 br_205 wl_106 vdd gnd cell_6t
Xbit_r107_c205 bl_205 br_205 wl_107 vdd gnd cell_6t
Xbit_r108_c205 bl_205 br_205 wl_108 vdd gnd cell_6t
Xbit_r109_c205 bl_205 br_205 wl_109 vdd gnd cell_6t
Xbit_r110_c205 bl_205 br_205 wl_110 vdd gnd cell_6t
Xbit_r111_c205 bl_205 br_205 wl_111 vdd gnd cell_6t
Xbit_r112_c205 bl_205 br_205 wl_112 vdd gnd cell_6t
Xbit_r113_c205 bl_205 br_205 wl_113 vdd gnd cell_6t
Xbit_r114_c205 bl_205 br_205 wl_114 vdd gnd cell_6t
Xbit_r115_c205 bl_205 br_205 wl_115 vdd gnd cell_6t
Xbit_r116_c205 bl_205 br_205 wl_116 vdd gnd cell_6t
Xbit_r117_c205 bl_205 br_205 wl_117 vdd gnd cell_6t
Xbit_r118_c205 bl_205 br_205 wl_118 vdd gnd cell_6t
Xbit_r119_c205 bl_205 br_205 wl_119 vdd gnd cell_6t
Xbit_r120_c205 bl_205 br_205 wl_120 vdd gnd cell_6t
Xbit_r121_c205 bl_205 br_205 wl_121 vdd gnd cell_6t
Xbit_r122_c205 bl_205 br_205 wl_122 vdd gnd cell_6t
Xbit_r123_c205 bl_205 br_205 wl_123 vdd gnd cell_6t
Xbit_r124_c205 bl_205 br_205 wl_124 vdd gnd cell_6t
Xbit_r125_c205 bl_205 br_205 wl_125 vdd gnd cell_6t
Xbit_r126_c205 bl_205 br_205 wl_126 vdd gnd cell_6t
Xbit_r127_c205 bl_205 br_205 wl_127 vdd gnd cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd cell_6t
Xbit_r1_c206 bl_206 br_206 wl_1 vdd gnd cell_6t
Xbit_r2_c206 bl_206 br_206 wl_2 vdd gnd cell_6t
Xbit_r3_c206 bl_206 br_206 wl_3 vdd gnd cell_6t
Xbit_r4_c206 bl_206 br_206 wl_4 vdd gnd cell_6t
Xbit_r5_c206 bl_206 br_206 wl_5 vdd gnd cell_6t
Xbit_r6_c206 bl_206 br_206 wl_6 vdd gnd cell_6t
Xbit_r7_c206 bl_206 br_206 wl_7 vdd gnd cell_6t
Xbit_r8_c206 bl_206 br_206 wl_8 vdd gnd cell_6t
Xbit_r9_c206 bl_206 br_206 wl_9 vdd gnd cell_6t
Xbit_r10_c206 bl_206 br_206 wl_10 vdd gnd cell_6t
Xbit_r11_c206 bl_206 br_206 wl_11 vdd gnd cell_6t
Xbit_r12_c206 bl_206 br_206 wl_12 vdd gnd cell_6t
Xbit_r13_c206 bl_206 br_206 wl_13 vdd gnd cell_6t
Xbit_r14_c206 bl_206 br_206 wl_14 vdd gnd cell_6t
Xbit_r15_c206 bl_206 br_206 wl_15 vdd gnd cell_6t
Xbit_r16_c206 bl_206 br_206 wl_16 vdd gnd cell_6t
Xbit_r17_c206 bl_206 br_206 wl_17 vdd gnd cell_6t
Xbit_r18_c206 bl_206 br_206 wl_18 vdd gnd cell_6t
Xbit_r19_c206 bl_206 br_206 wl_19 vdd gnd cell_6t
Xbit_r20_c206 bl_206 br_206 wl_20 vdd gnd cell_6t
Xbit_r21_c206 bl_206 br_206 wl_21 vdd gnd cell_6t
Xbit_r22_c206 bl_206 br_206 wl_22 vdd gnd cell_6t
Xbit_r23_c206 bl_206 br_206 wl_23 vdd gnd cell_6t
Xbit_r24_c206 bl_206 br_206 wl_24 vdd gnd cell_6t
Xbit_r25_c206 bl_206 br_206 wl_25 vdd gnd cell_6t
Xbit_r26_c206 bl_206 br_206 wl_26 vdd gnd cell_6t
Xbit_r27_c206 bl_206 br_206 wl_27 vdd gnd cell_6t
Xbit_r28_c206 bl_206 br_206 wl_28 vdd gnd cell_6t
Xbit_r29_c206 bl_206 br_206 wl_29 vdd gnd cell_6t
Xbit_r30_c206 bl_206 br_206 wl_30 vdd gnd cell_6t
Xbit_r31_c206 bl_206 br_206 wl_31 vdd gnd cell_6t
Xbit_r32_c206 bl_206 br_206 wl_32 vdd gnd cell_6t
Xbit_r33_c206 bl_206 br_206 wl_33 vdd gnd cell_6t
Xbit_r34_c206 bl_206 br_206 wl_34 vdd gnd cell_6t
Xbit_r35_c206 bl_206 br_206 wl_35 vdd gnd cell_6t
Xbit_r36_c206 bl_206 br_206 wl_36 vdd gnd cell_6t
Xbit_r37_c206 bl_206 br_206 wl_37 vdd gnd cell_6t
Xbit_r38_c206 bl_206 br_206 wl_38 vdd gnd cell_6t
Xbit_r39_c206 bl_206 br_206 wl_39 vdd gnd cell_6t
Xbit_r40_c206 bl_206 br_206 wl_40 vdd gnd cell_6t
Xbit_r41_c206 bl_206 br_206 wl_41 vdd gnd cell_6t
Xbit_r42_c206 bl_206 br_206 wl_42 vdd gnd cell_6t
Xbit_r43_c206 bl_206 br_206 wl_43 vdd gnd cell_6t
Xbit_r44_c206 bl_206 br_206 wl_44 vdd gnd cell_6t
Xbit_r45_c206 bl_206 br_206 wl_45 vdd gnd cell_6t
Xbit_r46_c206 bl_206 br_206 wl_46 vdd gnd cell_6t
Xbit_r47_c206 bl_206 br_206 wl_47 vdd gnd cell_6t
Xbit_r48_c206 bl_206 br_206 wl_48 vdd gnd cell_6t
Xbit_r49_c206 bl_206 br_206 wl_49 vdd gnd cell_6t
Xbit_r50_c206 bl_206 br_206 wl_50 vdd gnd cell_6t
Xbit_r51_c206 bl_206 br_206 wl_51 vdd gnd cell_6t
Xbit_r52_c206 bl_206 br_206 wl_52 vdd gnd cell_6t
Xbit_r53_c206 bl_206 br_206 wl_53 vdd gnd cell_6t
Xbit_r54_c206 bl_206 br_206 wl_54 vdd gnd cell_6t
Xbit_r55_c206 bl_206 br_206 wl_55 vdd gnd cell_6t
Xbit_r56_c206 bl_206 br_206 wl_56 vdd gnd cell_6t
Xbit_r57_c206 bl_206 br_206 wl_57 vdd gnd cell_6t
Xbit_r58_c206 bl_206 br_206 wl_58 vdd gnd cell_6t
Xbit_r59_c206 bl_206 br_206 wl_59 vdd gnd cell_6t
Xbit_r60_c206 bl_206 br_206 wl_60 vdd gnd cell_6t
Xbit_r61_c206 bl_206 br_206 wl_61 vdd gnd cell_6t
Xbit_r62_c206 bl_206 br_206 wl_62 vdd gnd cell_6t
Xbit_r63_c206 bl_206 br_206 wl_63 vdd gnd cell_6t
Xbit_r64_c206 bl_206 br_206 wl_64 vdd gnd cell_6t
Xbit_r65_c206 bl_206 br_206 wl_65 vdd gnd cell_6t
Xbit_r66_c206 bl_206 br_206 wl_66 vdd gnd cell_6t
Xbit_r67_c206 bl_206 br_206 wl_67 vdd gnd cell_6t
Xbit_r68_c206 bl_206 br_206 wl_68 vdd gnd cell_6t
Xbit_r69_c206 bl_206 br_206 wl_69 vdd gnd cell_6t
Xbit_r70_c206 bl_206 br_206 wl_70 vdd gnd cell_6t
Xbit_r71_c206 bl_206 br_206 wl_71 vdd gnd cell_6t
Xbit_r72_c206 bl_206 br_206 wl_72 vdd gnd cell_6t
Xbit_r73_c206 bl_206 br_206 wl_73 vdd gnd cell_6t
Xbit_r74_c206 bl_206 br_206 wl_74 vdd gnd cell_6t
Xbit_r75_c206 bl_206 br_206 wl_75 vdd gnd cell_6t
Xbit_r76_c206 bl_206 br_206 wl_76 vdd gnd cell_6t
Xbit_r77_c206 bl_206 br_206 wl_77 vdd gnd cell_6t
Xbit_r78_c206 bl_206 br_206 wl_78 vdd gnd cell_6t
Xbit_r79_c206 bl_206 br_206 wl_79 vdd gnd cell_6t
Xbit_r80_c206 bl_206 br_206 wl_80 vdd gnd cell_6t
Xbit_r81_c206 bl_206 br_206 wl_81 vdd gnd cell_6t
Xbit_r82_c206 bl_206 br_206 wl_82 vdd gnd cell_6t
Xbit_r83_c206 bl_206 br_206 wl_83 vdd gnd cell_6t
Xbit_r84_c206 bl_206 br_206 wl_84 vdd gnd cell_6t
Xbit_r85_c206 bl_206 br_206 wl_85 vdd gnd cell_6t
Xbit_r86_c206 bl_206 br_206 wl_86 vdd gnd cell_6t
Xbit_r87_c206 bl_206 br_206 wl_87 vdd gnd cell_6t
Xbit_r88_c206 bl_206 br_206 wl_88 vdd gnd cell_6t
Xbit_r89_c206 bl_206 br_206 wl_89 vdd gnd cell_6t
Xbit_r90_c206 bl_206 br_206 wl_90 vdd gnd cell_6t
Xbit_r91_c206 bl_206 br_206 wl_91 vdd gnd cell_6t
Xbit_r92_c206 bl_206 br_206 wl_92 vdd gnd cell_6t
Xbit_r93_c206 bl_206 br_206 wl_93 vdd gnd cell_6t
Xbit_r94_c206 bl_206 br_206 wl_94 vdd gnd cell_6t
Xbit_r95_c206 bl_206 br_206 wl_95 vdd gnd cell_6t
Xbit_r96_c206 bl_206 br_206 wl_96 vdd gnd cell_6t
Xbit_r97_c206 bl_206 br_206 wl_97 vdd gnd cell_6t
Xbit_r98_c206 bl_206 br_206 wl_98 vdd gnd cell_6t
Xbit_r99_c206 bl_206 br_206 wl_99 vdd gnd cell_6t
Xbit_r100_c206 bl_206 br_206 wl_100 vdd gnd cell_6t
Xbit_r101_c206 bl_206 br_206 wl_101 vdd gnd cell_6t
Xbit_r102_c206 bl_206 br_206 wl_102 vdd gnd cell_6t
Xbit_r103_c206 bl_206 br_206 wl_103 vdd gnd cell_6t
Xbit_r104_c206 bl_206 br_206 wl_104 vdd gnd cell_6t
Xbit_r105_c206 bl_206 br_206 wl_105 vdd gnd cell_6t
Xbit_r106_c206 bl_206 br_206 wl_106 vdd gnd cell_6t
Xbit_r107_c206 bl_206 br_206 wl_107 vdd gnd cell_6t
Xbit_r108_c206 bl_206 br_206 wl_108 vdd gnd cell_6t
Xbit_r109_c206 bl_206 br_206 wl_109 vdd gnd cell_6t
Xbit_r110_c206 bl_206 br_206 wl_110 vdd gnd cell_6t
Xbit_r111_c206 bl_206 br_206 wl_111 vdd gnd cell_6t
Xbit_r112_c206 bl_206 br_206 wl_112 vdd gnd cell_6t
Xbit_r113_c206 bl_206 br_206 wl_113 vdd gnd cell_6t
Xbit_r114_c206 bl_206 br_206 wl_114 vdd gnd cell_6t
Xbit_r115_c206 bl_206 br_206 wl_115 vdd gnd cell_6t
Xbit_r116_c206 bl_206 br_206 wl_116 vdd gnd cell_6t
Xbit_r117_c206 bl_206 br_206 wl_117 vdd gnd cell_6t
Xbit_r118_c206 bl_206 br_206 wl_118 vdd gnd cell_6t
Xbit_r119_c206 bl_206 br_206 wl_119 vdd gnd cell_6t
Xbit_r120_c206 bl_206 br_206 wl_120 vdd gnd cell_6t
Xbit_r121_c206 bl_206 br_206 wl_121 vdd gnd cell_6t
Xbit_r122_c206 bl_206 br_206 wl_122 vdd gnd cell_6t
Xbit_r123_c206 bl_206 br_206 wl_123 vdd gnd cell_6t
Xbit_r124_c206 bl_206 br_206 wl_124 vdd gnd cell_6t
Xbit_r125_c206 bl_206 br_206 wl_125 vdd gnd cell_6t
Xbit_r126_c206 bl_206 br_206 wl_126 vdd gnd cell_6t
Xbit_r127_c206 bl_206 br_206 wl_127 vdd gnd cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd cell_6t
Xbit_r1_c207 bl_207 br_207 wl_1 vdd gnd cell_6t
Xbit_r2_c207 bl_207 br_207 wl_2 vdd gnd cell_6t
Xbit_r3_c207 bl_207 br_207 wl_3 vdd gnd cell_6t
Xbit_r4_c207 bl_207 br_207 wl_4 vdd gnd cell_6t
Xbit_r5_c207 bl_207 br_207 wl_5 vdd gnd cell_6t
Xbit_r6_c207 bl_207 br_207 wl_6 vdd gnd cell_6t
Xbit_r7_c207 bl_207 br_207 wl_7 vdd gnd cell_6t
Xbit_r8_c207 bl_207 br_207 wl_8 vdd gnd cell_6t
Xbit_r9_c207 bl_207 br_207 wl_9 vdd gnd cell_6t
Xbit_r10_c207 bl_207 br_207 wl_10 vdd gnd cell_6t
Xbit_r11_c207 bl_207 br_207 wl_11 vdd gnd cell_6t
Xbit_r12_c207 bl_207 br_207 wl_12 vdd gnd cell_6t
Xbit_r13_c207 bl_207 br_207 wl_13 vdd gnd cell_6t
Xbit_r14_c207 bl_207 br_207 wl_14 vdd gnd cell_6t
Xbit_r15_c207 bl_207 br_207 wl_15 vdd gnd cell_6t
Xbit_r16_c207 bl_207 br_207 wl_16 vdd gnd cell_6t
Xbit_r17_c207 bl_207 br_207 wl_17 vdd gnd cell_6t
Xbit_r18_c207 bl_207 br_207 wl_18 vdd gnd cell_6t
Xbit_r19_c207 bl_207 br_207 wl_19 vdd gnd cell_6t
Xbit_r20_c207 bl_207 br_207 wl_20 vdd gnd cell_6t
Xbit_r21_c207 bl_207 br_207 wl_21 vdd gnd cell_6t
Xbit_r22_c207 bl_207 br_207 wl_22 vdd gnd cell_6t
Xbit_r23_c207 bl_207 br_207 wl_23 vdd gnd cell_6t
Xbit_r24_c207 bl_207 br_207 wl_24 vdd gnd cell_6t
Xbit_r25_c207 bl_207 br_207 wl_25 vdd gnd cell_6t
Xbit_r26_c207 bl_207 br_207 wl_26 vdd gnd cell_6t
Xbit_r27_c207 bl_207 br_207 wl_27 vdd gnd cell_6t
Xbit_r28_c207 bl_207 br_207 wl_28 vdd gnd cell_6t
Xbit_r29_c207 bl_207 br_207 wl_29 vdd gnd cell_6t
Xbit_r30_c207 bl_207 br_207 wl_30 vdd gnd cell_6t
Xbit_r31_c207 bl_207 br_207 wl_31 vdd gnd cell_6t
Xbit_r32_c207 bl_207 br_207 wl_32 vdd gnd cell_6t
Xbit_r33_c207 bl_207 br_207 wl_33 vdd gnd cell_6t
Xbit_r34_c207 bl_207 br_207 wl_34 vdd gnd cell_6t
Xbit_r35_c207 bl_207 br_207 wl_35 vdd gnd cell_6t
Xbit_r36_c207 bl_207 br_207 wl_36 vdd gnd cell_6t
Xbit_r37_c207 bl_207 br_207 wl_37 vdd gnd cell_6t
Xbit_r38_c207 bl_207 br_207 wl_38 vdd gnd cell_6t
Xbit_r39_c207 bl_207 br_207 wl_39 vdd gnd cell_6t
Xbit_r40_c207 bl_207 br_207 wl_40 vdd gnd cell_6t
Xbit_r41_c207 bl_207 br_207 wl_41 vdd gnd cell_6t
Xbit_r42_c207 bl_207 br_207 wl_42 vdd gnd cell_6t
Xbit_r43_c207 bl_207 br_207 wl_43 vdd gnd cell_6t
Xbit_r44_c207 bl_207 br_207 wl_44 vdd gnd cell_6t
Xbit_r45_c207 bl_207 br_207 wl_45 vdd gnd cell_6t
Xbit_r46_c207 bl_207 br_207 wl_46 vdd gnd cell_6t
Xbit_r47_c207 bl_207 br_207 wl_47 vdd gnd cell_6t
Xbit_r48_c207 bl_207 br_207 wl_48 vdd gnd cell_6t
Xbit_r49_c207 bl_207 br_207 wl_49 vdd gnd cell_6t
Xbit_r50_c207 bl_207 br_207 wl_50 vdd gnd cell_6t
Xbit_r51_c207 bl_207 br_207 wl_51 vdd gnd cell_6t
Xbit_r52_c207 bl_207 br_207 wl_52 vdd gnd cell_6t
Xbit_r53_c207 bl_207 br_207 wl_53 vdd gnd cell_6t
Xbit_r54_c207 bl_207 br_207 wl_54 vdd gnd cell_6t
Xbit_r55_c207 bl_207 br_207 wl_55 vdd gnd cell_6t
Xbit_r56_c207 bl_207 br_207 wl_56 vdd gnd cell_6t
Xbit_r57_c207 bl_207 br_207 wl_57 vdd gnd cell_6t
Xbit_r58_c207 bl_207 br_207 wl_58 vdd gnd cell_6t
Xbit_r59_c207 bl_207 br_207 wl_59 vdd gnd cell_6t
Xbit_r60_c207 bl_207 br_207 wl_60 vdd gnd cell_6t
Xbit_r61_c207 bl_207 br_207 wl_61 vdd gnd cell_6t
Xbit_r62_c207 bl_207 br_207 wl_62 vdd gnd cell_6t
Xbit_r63_c207 bl_207 br_207 wl_63 vdd gnd cell_6t
Xbit_r64_c207 bl_207 br_207 wl_64 vdd gnd cell_6t
Xbit_r65_c207 bl_207 br_207 wl_65 vdd gnd cell_6t
Xbit_r66_c207 bl_207 br_207 wl_66 vdd gnd cell_6t
Xbit_r67_c207 bl_207 br_207 wl_67 vdd gnd cell_6t
Xbit_r68_c207 bl_207 br_207 wl_68 vdd gnd cell_6t
Xbit_r69_c207 bl_207 br_207 wl_69 vdd gnd cell_6t
Xbit_r70_c207 bl_207 br_207 wl_70 vdd gnd cell_6t
Xbit_r71_c207 bl_207 br_207 wl_71 vdd gnd cell_6t
Xbit_r72_c207 bl_207 br_207 wl_72 vdd gnd cell_6t
Xbit_r73_c207 bl_207 br_207 wl_73 vdd gnd cell_6t
Xbit_r74_c207 bl_207 br_207 wl_74 vdd gnd cell_6t
Xbit_r75_c207 bl_207 br_207 wl_75 vdd gnd cell_6t
Xbit_r76_c207 bl_207 br_207 wl_76 vdd gnd cell_6t
Xbit_r77_c207 bl_207 br_207 wl_77 vdd gnd cell_6t
Xbit_r78_c207 bl_207 br_207 wl_78 vdd gnd cell_6t
Xbit_r79_c207 bl_207 br_207 wl_79 vdd gnd cell_6t
Xbit_r80_c207 bl_207 br_207 wl_80 vdd gnd cell_6t
Xbit_r81_c207 bl_207 br_207 wl_81 vdd gnd cell_6t
Xbit_r82_c207 bl_207 br_207 wl_82 vdd gnd cell_6t
Xbit_r83_c207 bl_207 br_207 wl_83 vdd gnd cell_6t
Xbit_r84_c207 bl_207 br_207 wl_84 vdd gnd cell_6t
Xbit_r85_c207 bl_207 br_207 wl_85 vdd gnd cell_6t
Xbit_r86_c207 bl_207 br_207 wl_86 vdd gnd cell_6t
Xbit_r87_c207 bl_207 br_207 wl_87 vdd gnd cell_6t
Xbit_r88_c207 bl_207 br_207 wl_88 vdd gnd cell_6t
Xbit_r89_c207 bl_207 br_207 wl_89 vdd gnd cell_6t
Xbit_r90_c207 bl_207 br_207 wl_90 vdd gnd cell_6t
Xbit_r91_c207 bl_207 br_207 wl_91 vdd gnd cell_6t
Xbit_r92_c207 bl_207 br_207 wl_92 vdd gnd cell_6t
Xbit_r93_c207 bl_207 br_207 wl_93 vdd gnd cell_6t
Xbit_r94_c207 bl_207 br_207 wl_94 vdd gnd cell_6t
Xbit_r95_c207 bl_207 br_207 wl_95 vdd gnd cell_6t
Xbit_r96_c207 bl_207 br_207 wl_96 vdd gnd cell_6t
Xbit_r97_c207 bl_207 br_207 wl_97 vdd gnd cell_6t
Xbit_r98_c207 bl_207 br_207 wl_98 vdd gnd cell_6t
Xbit_r99_c207 bl_207 br_207 wl_99 vdd gnd cell_6t
Xbit_r100_c207 bl_207 br_207 wl_100 vdd gnd cell_6t
Xbit_r101_c207 bl_207 br_207 wl_101 vdd gnd cell_6t
Xbit_r102_c207 bl_207 br_207 wl_102 vdd gnd cell_6t
Xbit_r103_c207 bl_207 br_207 wl_103 vdd gnd cell_6t
Xbit_r104_c207 bl_207 br_207 wl_104 vdd gnd cell_6t
Xbit_r105_c207 bl_207 br_207 wl_105 vdd gnd cell_6t
Xbit_r106_c207 bl_207 br_207 wl_106 vdd gnd cell_6t
Xbit_r107_c207 bl_207 br_207 wl_107 vdd gnd cell_6t
Xbit_r108_c207 bl_207 br_207 wl_108 vdd gnd cell_6t
Xbit_r109_c207 bl_207 br_207 wl_109 vdd gnd cell_6t
Xbit_r110_c207 bl_207 br_207 wl_110 vdd gnd cell_6t
Xbit_r111_c207 bl_207 br_207 wl_111 vdd gnd cell_6t
Xbit_r112_c207 bl_207 br_207 wl_112 vdd gnd cell_6t
Xbit_r113_c207 bl_207 br_207 wl_113 vdd gnd cell_6t
Xbit_r114_c207 bl_207 br_207 wl_114 vdd gnd cell_6t
Xbit_r115_c207 bl_207 br_207 wl_115 vdd gnd cell_6t
Xbit_r116_c207 bl_207 br_207 wl_116 vdd gnd cell_6t
Xbit_r117_c207 bl_207 br_207 wl_117 vdd gnd cell_6t
Xbit_r118_c207 bl_207 br_207 wl_118 vdd gnd cell_6t
Xbit_r119_c207 bl_207 br_207 wl_119 vdd gnd cell_6t
Xbit_r120_c207 bl_207 br_207 wl_120 vdd gnd cell_6t
Xbit_r121_c207 bl_207 br_207 wl_121 vdd gnd cell_6t
Xbit_r122_c207 bl_207 br_207 wl_122 vdd gnd cell_6t
Xbit_r123_c207 bl_207 br_207 wl_123 vdd gnd cell_6t
Xbit_r124_c207 bl_207 br_207 wl_124 vdd gnd cell_6t
Xbit_r125_c207 bl_207 br_207 wl_125 vdd gnd cell_6t
Xbit_r126_c207 bl_207 br_207 wl_126 vdd gnd cell_6t
Xbit_r127_c207 bl_207 br_207 wl_127 vdd gnd cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd cell_6t
Xbit_r1_c208 bl_208 br_208 wl_1 vdd gnd cell_6t
Xbit_r2_c208 bl_208 br_208 wl_2 vdd gnd cell_6t
Xbit_r3_c208 bl_208 br_208 wl_3 vdd gnd cell_6t
Xbit_r4_c208 bl_208 br_208 wl_4 vdd gnd cell_6t
Xbit_r5_c208 bl_208 br_208 wl_5 vdd gnd cell_6t
Xbit_r6_c208 bl_208 br_208 wl_6 vdd gnd cell_6t
Xbit_r7_c208 bl_208 br_208 wl_7 vdd gnd cell_6t
Xbit_r8_c208 bl_208 br_208 wl_8 vdd gnd cell_6t
Xbit_r9_c208 bl_208 br_208 wl_9 vdd gnd cell_6t
Xbit_r10_c208 bl_208 br_208 wl_10 vdd gnd cell_6t
Xbit_r11_c208 bl_208 br_208 wl_11 vdd gnd cell_6t
Xbit_r12_c208 bl_208 br_208 wl_12 vdd gnd cell_6t
Xbit_r13_c208 bl_208 br_208 wl_13 vdd gnd cell_6t
Xbit_r14_c208 bl_208 br_208 wl_14 vdd gnd cell_6t
Xbit_r15_c208 bl_208 br_208 wl_15 vdd gnd cell_6t
Xbit_r16_c208 bl_208 br_208 wl_16 vdd gnd cell_6t
Xbit_r17_c208 bl_208 br_208 wl_17 vdd gnd cell_6t
Xbit_r18_c208 bl_208 br_208 wl_18 vdd gnd cell_6t
Xbit_r19_c208 bl_208 br_208 wl_19 vdd gnd cell_6t
Xbit_r20_c208 bl_208 br_208 wl_20 vdd gnd cell_6t
Xbit_r21_c208 bl_208 br_208 wl_21 vdd gnd cell_6t
Xbit_r22_c208 bl_208 br_208 wl_22 vdd gnd cell_6t
Xbit_r23_c208 bl_208 br_208 wl_23 vdd gnd cell_6t
Xbit_r24_c208 bl_208 br_208 wl_24 vdd gnd cell_6t
Xbit_r25_c208 bl_208 br_208 wl_25 vdd gnd cell_6t
Xbit_r26_c208 bl_208 br_208 wl_26 vdd gnd cell_6t
Xbit_r27_c208 bl_208 br_208 wl_27 vdd gnd cell_6t
Xbit_r28_c208 bl_208 br_208 wl_28 vdd gnd cell_6t
Xbit_r29_c208 bl_208 br_208 wl_29 vdd gnd cell_6t
Xbit_r30_c208 bl_208 br_208 wl_30 vdd gnd cell_6t
Xbit_r31_c208 bl_208 br_208 wl_31 vdd gnd cell_6t
Xbit_r32_c208 bl_208 br_208 wl_32 vdd gnd cell_6t
Xbit_r33_c208 bl_208 br_208 wl_33 vdd gnd cell_6t
Xbit_r34_c208 bl_208 br_208 wl_34 vdd gnd cell_6t
Xbit_r35_c208 bl_208 br_208 wl_35 vdd gnd cell_6t
Xbit_r36_c208 bl_208 br_208 wl_36 vdd gnd cell_6t
Xbit_r37_c208 bl_208 br_208 wl_37 vdd gnd cell_6t
Xbit_r38_c208 bl_208 br_208 wl_38 vdd gnd cell_6t
Xbit_r39_c208 bl_208 br_208 wl_39 vdd gnd cell_6t
Xbit_r40_c208 bl_208 br_208 wl_40 vdd gnd cell_6t
Xbit_r41_c208 bl_208 br_208 wl_41 vdd gnd cell_6t
Xbit_r42_c208 bl_208 br_208 wl_42 vdd gnd cell_6t
Xbit_r43_c208 bl_208 br_208 wl_43 vdd gnd cell_6t
Xbit_r44_c208 bl_208 br_208 wl_44 vdd gnd cell_6t
Xbit_r45_c208 bl_208 br_208 wl_45 vdd gnd cell_6t
Xbit_r46_c208 bl_208 br_208 wl_46 vdd gnd cell_6t
Xbit_r47_c208 bl_208 br_208 wl_47 vdd gnd cell_6t
Xbit_r48_c208 bl_208 br_208 wl_48 vdd gnd cell_6t
Xbit_r49_c208 bl_208 br_208 wl_49 vdd gnd cell_6t
Xbit_r50_c208 bl_208 br_208 wl_50 vdd gnd cell_6t
Xbit_r51_c208 bl_208 br_208 wl_51 vdd gnd cell_6t
Xbit_r52_c208 bl_208 br_208 wl_52 vdd gnd cell_6t
Xbit_r53_c208 bl_208 br_208 wl_53 vdd gnd cell_6t
Xbit_r54_c208 bl_208 br_208 wl_54 vdd gnd cell_6t
Xbit_r55_c208 bl_208 br_208 wl_55 vdd gnd cell_6t
Xbit_r56_c208 bl_208 br_208 wl_56 vdd gnd cell_6t
Xbit_r57_c208 bl_208 br_208 wl_57 vdd gnd cell_6t
Xbit_r58_c208 bl_208 br_208 wl_58 vdd gnd cell_6t
Xbit_r59_c208 bl_208 br_208 wl_59 vdd gnd cell_6t
Xbit_r60_c208 bl_208 br_208 wl_60 vdd gnd cell_6t
Xbit_r61_c208 bl_208 br_208 wl_61 vdd gnd cell_6t
Xbit_r62_c208 bl_208 br_208 wl_62 vdd gnd cell_6t
Xbit_r63_c208 bl_208 br_208 wl_63 vdd gnd cell_6t
Xbit_r64_c208 bl_208 br_208 wl_64 vdd gnd cell_6t
Xbit_r65_c208 bl_208 br_208 wl_65 vdd gnd cell_6t
Xbit_r66_c208 bl_208 br_208 wl_66 vdd gnd cell_6t
Xbit_r67_c208 bl_208 br_208 wl_67 vdd gnd cell_6t
Xbit_r68_c208 bl_208 br_208 wl_68 vdd gnd cell_6t
Xbit_r69_c208 bl_208 br_208 wl_69 vdd gnd cell_6t
Xbit_r70_c208 bl_208 br_208 wl_70 vdd gnd cell_6t
Xbit_r71_c208 bl_208 br_208 wl_71 vdd gnd cell_6t
Xbit_r72_c208 bl_208 br_208 wl_72 vdd gnd cell_6t
Xbit_r73_c208 bl_208 br_208 wl_73 vdd gnd cell_6t
Xbit_r74_c208 bl_208 br_208 wl_74 vdd gnd cell_6t
Xbit_r75_c208 bl_208 br_208 wl_75 vdd gnd cell_6t
Xbit_r76_c208 bl_208 br_208 wl_76 vdd gnd cell_6t
Xbit_r77_c208 bl_208 br_208 wl_77 vdd gnd cell_6t
Xbit_r78_c208 bl_208 br_208 wl_78 vdd gnd cell_6t
Xbit_r79_c208 bl_208 br_208 wl_79 vdd gnd cell_6t
Xbit_r80_c208 bl_208 br_208 wl_80 vdd gnd cell_6t
Xbit_r81_c208 bl_208 br_208 wl_81 vdd gnd cell_6t
Xbit_r82_c208 bl_208 br_208 wl_82 vdd gnd cell_6t
Xbit_r83_c208 bl_208 br_208 wl_83 vdd gnd cell_6t
Xbit_r84_c208 bl_208 br_208 wl_84 vdd gnd cell_6t
Xbit_r85_c208 bl_208 br_208 wl_85 vdd gnd cell_6t
Xbit_r86_c208 bl_208 br_208 wl_86 vdd gnd cell_6t
Xbit_r87_c208 bl_208 br_208 wl_87 vdd gnd cell_6t
Xbit_r88_c208 bl_208 br_208 wl_88 vdd gnd cell_6t
Xbit_r89_c208 bl_208 br_208 wl_89 vdd gnd cell_6t
Xbit_r90_c208 bl_208 br_208 wl_90 vdd gnd cell_6t
Xbit_r91_c208 bl_208 br_208 wl_91 vdd gnd cell_6t
Xbit_r92_c208 bl_208 br_208 wl_92 vdd gnd cell_6t
Xbit_r93_c208 bl_208 br_208 wl_93 vdd gnd cell_6t
Xbit_r94_c208 bl_208 br_208 wl_94 vdd gnd cell_6t
Xbit_r95_c208 bl_208 br_208 wl_95 vdd gnd cell_6t
Xbit_r96_c208 bl_208 br_208 wl_96 vdd gnd cell_6t
Xbit_r97_c208 bl_208 br_208 wl_97 vdd gnd cell_6t
Xbit_r98_c208 bl_208 br_208 wl_98 vdd gnd cell_6t
Xbit_r99_c208 bl_208 br_208 wl_99 vdd gnd cell_6t
Xbit_r100_c208 bl_208 br_208 wl_100 vdd gnd cell_6t
Xbit_r101_c208 bl_208 br_208 wl_101 vdd gnd cell_6t
Xbit_r102_c208 bl_208 br_208 wl_102 vdd gnd cell_6t
Xbit_r103_c208 bl_208 br_208 wl_103 vdd gnd cell_6t
Xbit_r104_c208 bl_208 br_208 wl_104 vdd gnd cell_6t
Xbit_r105_c208 bl_208 br_208 wl_105 vdd gnd cell_6t
Xbit_r106_c208 bl_208 br_208 wl_106 vdd gnd cell_6t
Xbit_r107_c208 bl_208 br_208 wl_107 vdd gnd cell_6t
Xbit_r108_c208 bl_208 br_208 wl_108 vdd gnd cell_6t
Xbit_r109_c208 bl_208 br_208 wl_109 vdd gnd cell_6t
Xbit_r110_c208 bl_208 br_208 wl_110 vdd gnd cell_6t
Xbit_r111_c208 bl_208 br_208 wl_111 vdd gnd cell_6t
Xbit_r112_c208 bl_208 br_208 wl_112 vdd gnd cell_6t
Xbit_r113_c208 bl_208 br_208 wl_113 vdd gnd cell_6t
Xbit_r114_c208 bl_208 br_208 wl_114 vdd gnd cell_6t
Xbit_r115_c208 bl_208 br_208 wl_115 vdd gnd cell_6t
Xbit_r116_c208 bl_208 br_208 wl_116 vdd gnd cell_6t
Xbit_r117_c208 bl_208 br_208 wl_117 vdd gnd cell_6t
Xbit_r118_c208 bl_208 br_208 wl_118 vdd gnd cell_6t
Xbit_r119_c208 bl_208 br_208 wl_119 vdd gnd cell_6t
Xbit_r120_c208 bl_208 br_208 wl_120 vdd gnd cell_6t
Xbit_r121_c208 bl_208 br_208 wl_121 vdd gnd cell_6t
Xbit_r122_c208 bl_208 br_208 wl_122 vdd gnd cell_6t
Xbit_r123_c208 bl_208 br_208 wl_123 vdd gnd cell_6t
Xbit_r124_c208 bl_208 br_208 wl_124 vdd gnd cell_6t
Xbit_r125_c208 bl_208 br_208 wl_125 vdd gnd cell_6t
Xbit_r126_c208 bl_208 br_208 wl_126 vdd gnd cell_6t
Xbit_r127_c208 bl_208 br_208 wl_127 vdd gnd cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd cell_6t
Xbit_r1_c209 bl_209 br_209 wl_1 vdd gnd cell_6t
Xbit_r2_c209 bl_209 br_209 wl_2 vdd gnd cell_6t
Xbit_r3_c209 bl_209 br_209 wl_3 vdd gnd cell_6t
Xbit_r4_c209 bl_209 br_209 wl_4 vdd gnd cell_6t
Xbit_r5_c209 bl_209 br_209 wl_5 vdd gnd cell_6t
Xbit_r6_c209 bl_209 br_209 wl_6 vdd gnd cell_6t
Xbit_r7_c209 bl_209 br_209 wl_7 vdd gnd cell_6t
Xbit_r8_c209 bl_209 br_209 wl_8 vdd gnd cell_6t
Xbit_r9_c209 bl_209 br_209 wl_9 vdd gnd cell_6t
Xbit_r10_c209 bl_209 br_209 wl_10 vdd gnd cell_6t
Xbit_r11_c209 bl_209 br_209 wl_11 vdd gnd cell_6t
Xbit_r12_c209 bl_209 br_209 wl_12 vdd gnd cell_6t
Xbit_r13_c209 bl_209 br_209 wl_13 vdd gnd cell_6t
Xbit_r14_c209 bl_209 br_209 wl_14 vdd gnd cell_6t
Xbit_r15_c209 bl_209 br_209 wl_15 vdd gnd cell_6t
Xbit_r16_c209 bl_209 br_209 wl_16 vdd gnd cell_6t
Xbit_r17_c209 bl_209 br_209 wl_17 vdd gnd cell_6t
Xbit_r18_c209 bl_209 br_209 wl_18 vdd gnd cell_6t
Xbit_r19_c209 bl_209 br_209 wl_19 vdd gnd cell_6t
Xbit_r20_c209 bl_209 br_209 wl_20 vdd gnd cell_6t
Xbit_r21_c209 bl_209 br_209 wl_21 vdd gnd cell_6t
Xbit_r22_c209 bl_209 br_209 wl_22 vdd gnd cell_6t
Xbit_r23_c209 bl_209 br_209 wl_23 vdd gnd cell_6t
Xbit_r24_c209 bl_209 br_209 wl_24 vdd gnd cell_6t
Xbit_r25_c209 bl_209 br_209 wl_25 vdd gnd cell_6t
Xbit_r26_c209 bl_209 br_209 wl_26 vdd gnd cell_6t
Xbit_r27_c209 bl_209 br_209 wl_27 vdd gnd cell_6t
Xbit_r28_c209 bl_209 br_209 wl_28 vdd gnd cell_6t
Xbit_r29_c209 bl_209 br_209 wl_29 vdd gnd cell_6t
Xbit_r30_c209 bl_209 br_209 wl_30 vdd gnd cell_6t
Xbit_r31_c209 bl_209 br_209 wl_31 vdd gnd cell_6t
Xbit_r32_c209 bl_209 br_209 wl_32 vdd gnd cell_6t
Xbit_r33_c209 bl_209 br_209 wl_33 vdd gnd cell_6t
Xbit_r34_c209 bl_209 br_209 wl_34 vdd gnd cell_6t
Xbit_r35_c209 bl_209 br_209 wl_35 vdd gnd cell_6t
Xbit_r36_c209 bl_209 br_209 wl_36 vdd gnd cell_6t
Xbit_r37_c209 bl_209 br_209 wl_37 vdd gnd cell_6t
Xbit_r38_c209 bl_209 br_209 wl_38 vdd gnd cell_6t
Xbit_r39_c209 bl_209 br_209 wl_39 vdd gnd cell_6t
Xbit_r40_c209 bl_209 br_209 wl_40 vdd gnd cell_6t
Xbit_r41_c209 bl_209 br_209 wl_41 vdd gnd cell_6t
Xbit_r42_c209 bl_209 br_209 wl_42 vdd gnd cell_6t
Xbit_r43_c209 bl_209 br_209 wl_43 vdd gnd cell_6t
Xbit_r44_c209 bl_209 br_209 wl_44 vdd gnd cell_6t
Xbit_r45_c209 bl_209 br_209 wl_45 vdd gnd cell_6t
Xbit_r46_c209 bl_209 br_209 wl_46 vdd gnd cell_6t
Xbit_r47_c209 bl_209 br_209 wl_47 vdd gnd cell_6t
Xbit_r48_c209 bl_209 br_209 wl_48 vdd gnd cell_6t
Xbit_r49_c209 bl_209 br_209 wl_49 vdd gnd cell_6t
Xbit_r50_c209 bl_209 br_209 wl_50 vdd gnd cell_6t
Xbit_r51_c209 bl_209 br_209 wl_51 vdd gnd cell_6t
Xbit_r52_c209 bl_209 br_209 wl_52 vdd gnd cell_6t
Xbit_r53_c209 bl_209 br_209 wl_53 vdd gnd cell_6t
Xbit_r54_c209 bl_209 br_209 wl_54 vdd gnd cell_6t
Xbit_r55_c209 bl_209 br_209 wl_55 vdd gnd cell_6t
Xbit_r56_c209 bl_209 br_209 wl_56 vdd gnd cell_6t
Xbit_r57_c209 bl_209 br_209 wl_57 vdd gnd cell_6t
Xbit_r58_c209 bl_209 br_209 wl_58 vdd gnd cell_6t
Xbit_r59_c209 bl_209 br_209 wl_59 vdd gnd cell_6t
Xbit_r60_c209 bl_209 br_209 wl_60 vdd gnd cell_6t
Xbit_r61_c209 bl_209 br_209 wl_61 vdd gnd cell_6t
Xbit_r62_c209 bl_209 br_209 wl_62 vdd gnd cell_6t
Xbit_r63_c209 bl_209 br_209 wl_63 vdd gnd cell_6t
Xbit_r64_c209 bl_209 br_209 wl_64 vdd gnd cell_6t
Xbit_r65_c209 bl_209 br_209 wl_65 vdd gnd cell_6t
Xbit_r66_c209 bl_209 br_209 wl_66 vdd gnd cell_6t
Xbit_r67_c209 bl_209 br_209 wl_67 vdd gnd cell_6t
Xbit_r68_c209 bl_209 br_209 wl_68 vdd gnd cell_6t
Xbit_r69_c209 bl_209 br_209 wl_69 vdd gnd cell_6t
Xbit_r70_c209 bl_209 br_209 wl_70 vdd gnd cell_6t
Xbit_r71_c209 bl_209 br_209 wl_71 vdd gnd cell_6t
Xbit_r72_c209 bl_209 br_209 wl_72 vdd gnd cell_6t
Xbit_r73_c209 bl_209 br_209 wl_73 vdd gnd cell_6t
Xbit_r74_c209 bl_209 br_209 wl_74 vdd gnd cell_6t
Xbit_r75_c209 bl_209 br_209 wl_75 vdd gnd cell_6t
Xbit_r76_c209 bl_209 br_209 wl_76 vdd gnd cell_6t
Xbit_r77_c209 bl_209 br_209 wl_77 vdd gnd cell_6t
Xbit_r78_c209 bl_209 br_209 wl_78 vdd gnd cell_6t
Xbit_r79_c209 bl_209 br_209 wl_79 vdd gnd cell_6t
Xbit_r80_c209 bl_209 br_209 wl_80 vdd gnd cell_6t
Xbit_r81_c209 bl_209 br_209 wl_81 vdd gnd cell_6t
Xbit_r82_c209 bl_209 br_209 wl_82 vdd gnd cell_6t
Xbit_r83_c209 bl_209 br_209 wl_83 vdd gnd cell_6t
Xbit_r84_c209 bl_209 br_209 wl_84 vdd gnd cell_6t
Xbit_r85_c209 bl_209 br_209 wl_85 vdd gnd cell_6t
Xbit_r86_c209 bl_209 br_209 wl_86 vdd gnd cell_6t
Xbit_r87_c209 bl_209 br_209 wl_87 vdd gnd cell_6t
Xbit_r88_c209 bl_209 br_209 wl_88 vdd gnd cell_6t
Xbit_r89_c209 bl_209 br_209 wl_89 vdd gnd cell_6t
Xbit_r90_c209 bl_209 br_209 wl_90 vdd gnd cell_6t
Xbit_r91_c209 bl_209 br_209 wl_91 vdd gnd cell_6t
Xbit_r92_c209 bl_209 br_209 wl_92 vdd gnd cell_6t
Xbit_r93_c209 bl_209 br_209 wl_93 vdd gnd cell_6t
Xbit_r94_c209 bl_209 br_209 wl_94 vdd gnd cell_6t
Xbit_r95_c209 bl_209 br_209 wl_95 vdd gnd cell_6t
Xbit_r96_c209 bl_209 br_209 wl_96 vdd gnd cell_6t
Xbit_r97_c209 bl_209 br_209 wl_97 vdd gnd cell_6t
Xbit_r98_c209 bl_209 br_209 wl_98 vdd gnd cell_6t
Xbit_r99_c209 bl_209 br_209 wl_99 vdd gnd cell_6t
Xbit_r100_c209 bl_209 br_209 wl_100 vdd gnd cell_6t
Xbit_r101_c209 bl_209 br_209 wl_101 vdd gnd cell_6t
Xbit_r102_c209 bl_209 br_209 wl_102 vdd gnd cell_6t
Xbit_r103_c209 bl_209 br_209 wl_103 vdd gnd cell_6t
Xbit_r104_c209 bl_209 br_209 wl_104 vdd gnd cell_6t
Xbit_r105_c209 bl_209 br_209 wl_105 vdd gnd cell_6t
Xbit_r106_c209 bl_209 br_209 wl_106 vdd gnd cell_6t
Xbit_r107_c209 bl_209 br_209 wl_107 vdd gnd cell_6t
Xbit_r108_c209 bl_209 br_209 wl_108 vdd gnd cell_6t
Xbit_r109_c209 bl_209 br_209 wl_109 vdd gnd cell_6t
Xbit_r110_c209 bl_209 br_209 wl_110 vdd gnd cell_6t
Xbit_r111_c209 bl_209 br_209 wl_111 vdd gnd cell_6t
Xbit_r112_c209 bl_209 br_209 wl_112 vdd gnd cell_6t
Xbit_r113_c209 bl_209 br_209 wl_113 vdd gnd cell_6t
Xbit_r114_c209 bl_209 br_209 wl_114 vdd gnd cell_6t
Xbit_r115_c209 bl_209 br_209 wl_115 vdd gnd cell_6t
Xbit_r116_c209 bl_209 br_209 wl_116 vdd gnd cell_6t
Xbit_r117_c209 bl_209 br_209 wl_117 vdd gnd cell_6t
Xbit_r118_c209 bl_209 br_209 wl_118 vdd gnd cell_6t
Xbit_r119_c209 bl_209 br_209 wl_119 vdd gnd cell_6t
Xbit_r120_c209 bl_209 br_209 wl_120 vdd gnd cell_6t
Xbit_r121_c209 bl_209 br_209 wl_121 vdd gnd cell_6t
Xbit_r122_c209 bl_209 br_209 wl_122 vdd gnd cell_6t
Xbit_r123_c209 bl_209 br_209 wl_123 vdd gnd cell_6t
Xbit_r124_c209 bl_209 br_209 wl_124 vdd gnd cell_6t
Xbit_r125_c209 bl_209 br_209 wl_125 vdd gnd cell_6t
Xbit_r126_c209 bl_209 br_209 wl_126 vdd gnd cell_6t
Xbit_r127_c209 bl_209 br_209 wl_127 vdd gnd cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd cell_6t
Xbit_r1_c210 bl_210 br_210 wl_1 vdd gnd cell_6t
Xbit_r2_c210 bl_210 br_210 wl_2 vdd gnd cell_6t
Xbit_r3_c210 bl_210 br_210 wl_3 vdd gnd cell_6t
Xbit_r4_c210 bl_210 br_210 wl_4 vdd gnd cell_6t
Xbit_r5_c210 bl_210 br_210 wl_5 vdd gnd cell_6t
Xbit_r6_c210 bl_210 br_210 wl_6 vdd gnd cell_6t
Xbit_r7_c210 bl_210 br_210 wl_7 vdd gnd cell_6t
Xbit_r8_c210 bl_210 br_210 wl_8 vdd gnd cell_6t
Xbit_r9_c210 bl_210 br_210 wl_9 vdd gnd cell_6t
Xbit_r10_c210 bl_210 br_210 wl_10 vdd gnd cell_6t
Xbit_r11_c210 bl_210 br_210 wl_11 vdd gnd cell_6t
Xbit_r12_c210 bl_210 br_210 wl_12 vdd gnd cell_6t
Xbit_r13_c210 bl_210 br_210 wl_13 vdd gnd cell_6t
Xbit_r14_c210 bl_210 br_210 wl_14 vdd gnd cell_6t
Xbit_r15_c210 bl_210 br_210 wl_15 vdd gnd cell_6t
Xbit_r16_c210 bl_210 br_210 wl_16 vdd gnd cell_6t
Xbit_r17_c210 bl_210 br_210 wl_17 vdd gnd cell_6t
Xbit_r18_c210 bl_210 br_210 wl_18 vdd gnd cell_6t
Xbit_r19_c210 bl_210 br_210 wl_19 vdd gnd cell_6t
Xbit_r20_c210 bl_210 br_210 wl_20 vdd gnd cell_6t
Xbit_r21_c210 bl_210 br_210 wl_21 vdd gnd cell_6t
Xbit_r22_c210 bl_210 br_210 wl_22 vdd gnd cell_6t
Xbit_r23_c210 bl_210 br_210 wl_23 vdd gnd cell_6t
Xbit_r24_c210 bl_210 br_210 wl_24 vdd gnd cell_6t
Xbit_r25_c210 bl_210 br_210 wl_25 vdd gnd cell_6t
Xbit_r26_c210 bl_210 br_210 wl_26 vdd gnd cell_6t
Xbit_r27_c210 bl_210 br_210 wl_27 vdd gnd cell_6t
Xbit_r28_c210 bl_210 br_210 wl_28 vdd gnd cell_6t
Xbit_r29_c210 bl_210 br_210 wl_29 vdd gnd cell_6t
Xbit_r30_c210 bl_210 br_210 wl_30 vdd gnd cell_6t
Xbit_r31_c210 bl_210 br_210 wl_31 vdd gnd cell_6t
Xbit_r32_c210 bl_210 br_210 wl_32 vdd gnd cell_6t
Xbit_r33_c210 bl_210 br_210 wl_33 vdd gnd cell_6t
Xbit_r34_c210 bl_210 br_210 wl_34 vdd gnd cell_6t
Xbit_r35_c210 bl_210 br_210 wl_35 vdd gnd cell_6t
Xbit_r36_c210 bl_210 br_210 wl_36 vdd gnd cell_6t
Xbit_r37_c210 bl_210 br_210 wl_37 vdd gnd cell_6t
Xbit_r38_c210 bl_210 br_210 wl_38 vdd gnd cell_6t
Xbit_r39_c210 bl_210 br_210 wl_39 vdd gnd cell_6t
Xbit_r40_c210 bl_210 br_210 wl_40 vdd gnd cell_6t
Xbit_r41_c210 bl_210 br_210 wl_41 vdd gnd cell_6t
Xbit_r42_c210 bl_210 br_210 wl_42 vdd gnd cell_6t
Xbit_r43_c210 bl_210 br_210 wl_43 vdd gnd cell_6t
Xbit_r44_c210 bl_210 br_210 wl_44 vdd gnd cell_6t
Xbit_r45_c210 bl_210 br_210 wl_45 vdd gnd cell_6t
Xbit_r46_c210 bl_210 br_210 wl_46 vdd gnd cell_6t
Xbit_r47_c210 bl_210 br_210 wl_47 vdd gnd cell_6t
Xbit_r48_c210 bl_210 br_210 wl_48 vdd gnd cell_6t
Xbit_r49_c210 bl_210 br_210 wl_49 vdd gnd cell_6t
Xbit_r50_c210 bl_210 br_210 wl_50 vdd gnd cell_6t
Xbit_r51_c210 bl_210 br_210 wl_51 vdd gnd cell_6t
Xbit_r52_c210 bl_210 br_210 wl_52 vdd gnd cell_6t
Xbit_r53_c210 bl_210 br_210 wl_53 vdd gnd cell_6t
Xbit_r54_c210 bl_210 br_210 wl_54 vdd gnd cell_6t
Xbit_r55_c210 bl_210 br_210 wl_55 vdd gnd cell_6t
Xbit_r56_c210 bl_210 br_210 wl_56 vdd gnd cell_6t
Xbit_r57_c210 bl_210 br_210 wl_57 vdd gnd cell_6t
Xbit_r58_c210 bl_210 br_210 wl_58 vdd gnd cell_6t
Xbit_r59_c210 bl_210 br_210 wl_59 vdd gnd cell_6t
Xbit_r60_c210 bl_210 br_210 wl_60 vdd gnd cell_6t
Xbit_r61_c210 bl_210 br_210 wl_61 vdd gnd cell_6t
Xbit_r62_c210 bl_210 br_210 wl_62 vdd gnd cell_6t
Xbit_r63_c210 bl_210 br_210 wl_63 vdd gnd cell_6t
Xbit_r64_c210 bl_210 br_210 wl_64 vdd gnd cell_6t
Xbit_r65_c210 bl_210 br_210 wl_65 vdd gnd cell_6t
Xbit_r66_c210 bl_210 br_210 wl_66 vdd gnd cell_6t
Xbit_r67_c210 bl_210 br_210 wl_67 vdd gnd cell_6t
Xbit_r68_c210 bl_210 br_210 wl_68 vdd gnd cell_6t
Xbit_r69_c210 bl_210 br_210 wl_69 vdd gnd cell_6t
Xbit_r70_c210 bl_210 br_210 wl_70 vdd gnd cell_6t
Xbit_r71_c210 bl_210 br_210 wl_71 vdd gnd cell_6t
Xbit_r72_c210 bl_210 br_210 wl_72 vdd gnd cell_6t
Xbit_r73_c210 bl_210 br_210 wl_73 vdd gnd cell_6t
Xbit_r74_c210 bl_210 br_210 wl_74 vdd gnd cell_6t
Xbit_r75_c210 bl_210 br_210 wl_75 vdd gnd cell_6t
Xbit_r76_c210 bl_210 br_210 wl_76 vdd gnd cell_6t
Xbit_r77_c210 bl_210 br_210 wl_77 vdd gnd cell_6t
Xbit_r78_c210 bl_210 br_210 wl_78 vdd gnd cell_6t
Xbit_r79_c210 bl_210 br_210 wl_79 vdd gnd cell_6t
Xbit_r80_c210 bl_210 br_210 wl_80 vdd gnd cell_6t
Xbit_r81_c210 bl_210 br_210 wl_81 vdd gnd cell_6t
Xbit_r82_c210 bl_210 br_210 wl_82 vdd gnd cell_6t
Xbit_r83_c210 bl_210 br_210 wl_83 vdd gnd cell_6t
Xbit_r84_c210 bl_210 br_210 wl_84 vdd gnd cell_6t
Xbit_r85_c210 bl_210 br_210 wl_85 vdd gnd cell_6t
Xbit_r86_c210 bl_210 br_210 wl_86 vdd gnd cell_6t
Xbit_r87_c210 bl_210 br_210 wl_87 vdd gnd cell_6t
Xbit_r88_c210 bl_210 br_210 wl_88 vdd gnd cell_6t
Xbit_r89_c210 bl_210 br_210 wl_89 vdd gnd cell_6t
Xbit_r90_c210 bl_210 br_210 wl_90 vdd gnd cell_6t
Xbit_r91_c210 bl_210 br_210 wl_91 vdd gnd cell_6t
Xbit_r92_c210 bl_210 br_210 wl_92 vdd gnd cell_6t
Xbit_r93_c210 bl_210 br_210 wl_93 vdd gnd cell_6t
Xbit_r94_c210 bl_210 br_210 wl_94 vdd gnd cell_6t
Xbit_r95_c210 bl_210 br_210 wl_95 vdd gnd cell_6t
Xbit_r96_c210 bl_210 br_210 wl_96 vdd gnd cell_6t
Xbit_r97_c210 bl_210 br_210 wl_97 vdd gnd cell_6t
Xbit_r98_c210 bl_210 br_210 wl_98 vdd gnd cell_6t
Xbit_r99_c210 bl_210 br_210 wl_99 vdd gnd cell_6t
Xbit_r100_c210 bl_210 br_210 wl_100 vdd gnd cell_6t
Xbit_r101_c210 bl_210 br_210 wl_101 vdd gnd cell_6t
Xbit_r102_c210 bl_210 br_210 wl_102 vdd gnd cell_6t
Xbit_r103_c210 bl_210 br_210 wl_103 vdd gnd cell_6t
Xbit_r104_c210 bl_210 br_210 wl_104 vdd gnd cell_6t
Xbit_r105_c210 bl_210 br_210 wl_105 vdd gnd cell_6t
Xbit_r106_c210 bl_210 br_210 wl_106 vdd gnd cell_6t
Xbit_r107_c210 bl_210 br_210 wl_107 vdd gnd cell_6t
Xbit_r108_c210 bl_210 br_210 wl_108 vdd gnd cell_6t
Xbit_r109_c210 bl_210 br_210 wl_109 vdd gnd cell_6t
Xbit_r110_c210 bl_210 br_210 wl_110 vdd gnd cell_6t
Xbit_r111_c210 bl_210 br_210 wl_111 vdd gnd cell_6t
Xbit_r112_c210 bl_210 br_210 wl_112 vdd gnd cell_6t
Xbit_r113_c210 bl_210 br_210 wl_113 vdd gnd cell_6t
Xbit_r114_c210 bl_210 br_210 wl_114 vdd gnd cell_6t
Xbit_r115_c210 bl_210 br_210 wl_115 vdd gnd cell_6t
Xbit_r116_c210 bl_210 br_210 wl_116 vdd gnd cell_6t
Xbit_r117_c210 bl_210 br_210 wl_117 vdd gnd cell_6t
Xbit_r118_c210 bl_210 br_210 wl_118 vdd gnd cell_6t
Xbit_r119_c210 bl_210 br_210 wl_119 vdd gnd cell_6t
Xbit_r120_c210 bl_210 br_210 wl_120 vdd gnd cell_6t
Xbit_r121_c210 bl_210 br_210 wl_121 vdd gnd cell_6t
Xbit_r122_c210 bl_210 br_210 wl_122 vdd gnd cell_6t
Xbit_r123_c210 bl_210 br_210 wl_123 vdd gnd cell_6t
Xbit_r124_c210 bl_210 br_210 wl_124 vdd gnd cell_6t
Xbit_r125_c210 bl_210 br_210 wl_125 vdd gnd cell_6t
Xbit_r126_c210 bl_210 br_210 wl_126 vdd gnd cell_6t
Xbit_r127_c210 bl_210 br_210 wl_127 vdd gnd cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd cell_6t
Xbit_r1_c211 bl_211 br_211 wl_1 vdd gnd cell_6t
Xbit_r2_c211 bl_211 br_211 wl_2 vdd gnd cell_6t
Xbit_r3_c211 bl_211 br_211 wl_3 vdd gnd cell_6t
Xbit_r4_c211 bl_211 br_211 wl_4 vdd gnd cell_6t
Xbit_r5_c211 bl_211 br_211 wl_5 vdd gnd cell_6t
Xbit_r6_c211 bl_211 br_211 wl_6 vdd gnd cell_6t
Xbit_r7_c211 bl_211 br_211 wl_7 vdd gnd cell_6t
Xbit_r8_c211 bl_211 br_211 wl_8 vdd gnd cell_6t
Xbit_r9_c211 bl_211 br_211 wl_9 vdd gnd cell_6t
Xbit_r10_c211 bl_211 br_211 wl_10 vdd gnd cell_6t
Xbit_r11_c211 bl_211 br_211 wl_11 vdd gnd cell_6t
Xbit_r12_c211 bl_211 br_211 wl_12 vdd gnd cell_6t
Xbit_r13_c211 bl_211 br_211 wl_13 vdd gnd cell_6t
Xbit_r14_c211 bl_211 br_211 wl_14 vdd gnd cell_6t
Xbit_r15_c211 bl_211 br_211 wl_15 vdd gnd cell_6t
Xbit_r16_c211 bl_211 br_211 wl_16 vdd gnd cell_6t
Xbit_r17_c211 bl_211 br_211 wl_17 vdd gnd cell_6t
Xbit_r18_c211 bl_211 br_211 wl_18 vdd gnd cell_6t
Xbit_r19_c211 bl_211 br_211 wl_19 vdd gnd cell_6t
Xbit_r20_c211 bl_211 br_211 wl_20 vdd gnd cell_6t
Xbit_r21_c211 bl_211 br_211 wl_21 vdd gnd cell_6t
Xbit_r22_c211 bl_211 br_211 wl_22 vdd gnd cell_6t
Xbit_r23_c211 bl_211 br_211 wl_23 vdd gnd cell_6t
Xbit_r24_c211 bl_211 br_211 wl_24 vdd gnd cell_6t
Xbit_r25_c211 bl_211 br_211 wl_25 vdd gnd cell_6t
Xbit_r26_c211 bl_211 br_211 wl_26 vdd gnd cell_6t
Xbit_r27_c211 bl_211 br_211 wl_27 vdd gnd cell_6t
Xbit_r28_c211 bl_211 br_211 wl_28 vdd gnd cell_6t
Xbit_r29_c211 bl_211 br_211 wl_29 vdd gnd cell_6t
Xbit_r30_c211 bl_211 br_211 wl_30 vdd gnd cell_6t
Xbit_r31_c211 bl_211 br_211 wl_31 vdd gnd cell_6t
Xbit_r32_c211 bl_211 br_211 wl_32 vdd gnd cell_6t
Xbit_r33_c211 bl_211 br_211 wl_33 vdd gnd cell_6t
Xbit_r34_c211 bl_211 br_211 wl_34 vdd gnd cell_6t
Xbit_r35_c211 bl_211 br_211 wl_35 vdd gnd cell_6t
Xbit_r36_c211 bl_211 br_211 wl_36 vdd gnd cell_6t
Xbit_r37_c211 bl_211 br_211 wl_37 vdd gnd cell_6t
Xbit_r38_c211 bl_211 br_211 wl_38 vdd gnd cell_6t
Xbit_r39_c211 bl_211 br_211 wl_39 vdd gnd cell_6t
Xbit_r40_c211 bl_211 br_211 wl_40 vdd gnd cell_6t
Xbit_r41_c211 bl_211 br_211 wl_41 vdd gnd cell_6t
Xbit_r42_c211 bl_211 br_211 wl_42 vdd gnd cell_6t
Xbit_r43_c211 bl_211 br_211 wl_43 vdd gnd cell_6t
Xbit_r44_c211 bl_211 br_211 wl_44 vdd gnd cell_6t
Xbit_r45_c211 bl_211 br_211 wl_45 vdd gnd cell_6t
Xbit_r46_c211 bl_211 br_211 wl_46 vdd gnd cell_6t
Xbit_r47_c211 bl_211 br_211 wl_47 vdd gnd cell_6t
Xbit_r48_c211 bl_211 br_211 wl_48 vdd gnd cell_6t
Xbit_r49_c211 bl_211 br_211 wl_49 vdd gnd cell_6t
Xbit_r50_c211 bl_211 br_211 wl_50 vdd gnd cell_6t
Xbit_r51_c211 bl_211 br_211 wl_51 vdd gnd cell_6t
Xbit_r52_c211 bl_211 br_211 wl_52 vdd gnd cell_6t
Xbit_r53_c211 bl_211 br_211 wl_53 vdd gnd cell_6t
Xbit_r54_c211 bl_211 br_211 wl_54 vdd gnd cell_6t
Xbit_r55_c211 bl_211 br_211 wl_55 vdd gnd cell_6t
Xbit_r56_c211 bl_211 br_211 wl_56 vdd gnd cell_6t
Xbit_r57_c211 bl_211 br_211 wl_57 vdd gnd cell_6t
Xbit_r58_c211 bl_211 br_211 wl_58 vdd gnd cell_6t
Xbit_r59_c211 bl_211 br_211 wl_59 vdd gnd cell_6t
Xbit_r60_c211 bl_211 br_211 wl_60 vdd gnd cell_6t
Xbit_r61_c211 bl_211 br_211 wl_61 vdd gnd cell_6t
Xbit_r62_c211 bl_211 br_211 wl_62 vdd gnd cell_6t
Xbit_r63_c211 bl_211 br_211 wl_63 vdd gnd cell_6t
Xbit_r64_c211 bl_211 br_211 wl_64 vdd gnd cell_6t
Xbit_r65_c211 bl_211 br_211 wl_65 vdd gnd cell_6t
Xbit_r66_c211 bl_211 br_211 wl_66 vdd gnd cell_6t
Xbit_r67_c211 bl_211 br_211 wl_67 vdd gnd cell_6t
Xbit_r68_c211 bl_211 br_211 wl_68 vdd gnd cell_6t
Xbit_r69_c211 bl_211 br_211 wl_69 vdd gnd cell_6t
Xbit_r70_c211 bl_211 br_211 wl_70 vdd gnd cell_6t
Xbit_r71_c211 bl_211 br_211 wl_71 vdd gnd cell_6t
Xbit_r72_c211 bl_211 br_211 wl_72 vdd gnd cell_6t
Xbit_r73_c211 bl_211 br_211 wl_73 vdd gnd cell_6t
Xbit_r74_c211 bl_211 br_211 wl_74 vdd gnd cell_6t
Xbit_r75_c211 bl_211 br_211 wl_75 vdd gnd cell_6t
Xbit_r76_c211 bl_211 br_211 wl_76 vdd gnd cell_6t
Xbit_r77_c211 bl_211 br_211 wl_77 vdd gnd cell_6t
Xbit_r78_c211 bl_211 br_211 wl_78 vdd gnd cell_6t
Xbit_r79_c211 bl_211 br_211 wl_79 vdd gnd cell_6t
Xbit_r80_c211 bl_211 br_211 wl_80 vdd gnd cell_6t
Xbit_r81_c211 bl_211 br_211 wl_81 vdd gnd cell_6t
Xbit_r82_c211 bl_211 br_211 wl_82 vdd gnd cell_6t
Xbit_r83_c211 bl_211 br_211 wl_83 vdd gnd cell_6t
Xbit_r84_c211 bl_211 br_211 wl_84 vdd gnd cell_6t
Xbit_r85_c211 bl_211 br_211 wl_85 vdd gnd cell_6t
Xbit_r86_c211 bl_211 br_211 wl_86 vdd gnd cell_6t
Xbit_r87_c211 bl_211 br_211 wl_87 vdd gnd cell_6t
Xbit_r88_c211 bl_211 br_211 wl_88 vdd gnd cell_6t
Xbit_r89_c211 bl_211 br_211 wl_89 vdd gnd cell_6t
Xbit_r90_c211 bl_211 br_211 wl_90 vdd gnd cell_6t
Xbit_r91_c211 bl_211 br_211 wl_91 vdd gnd cell_6t
Xbit_r92_c211 bl_211 br_211 wl_92 vdd gnd cell_6t
Xbit_r93_c211 bl_211 br_211 wl_93 vdd gnd cell_6t
Xbit_r94_c211 bl_211 br_211 wl_94 vdd gnd cell_6t
Xbit_r95_c211 bl_211 br_211 wl_95 vdd gnd cell_6t
Xbit_r96_c211 bl_211 br_211 wl_96 vdd gnd cell_6t
Xbit_r97_c211 bl_211 br_211 wl_97 vdd gnd cell_6t
Xbit_r98_c211 bl_211 br_211 wl_98 vdd gnd cell_6t
Xbit_r99_c211 bl_211 br_211 wl_99 vdd gnd cell_6t
Xbit_r100_c211 bl_211 br_211 wl_100 vdd gnd cell_6t
Xbit_r101_c211 bl_211 br_211 wl_101 vdd gnd cell_6t
Xbit_r102_c211 bl_211 br_211 wl_102 vdd gnd cell_6t
Xbit_r103_c211 bl_211 br_211 wl_103 vdd gnd cell_6t
Xbit_r104_c211 bl_211 br_211 wl_104 vdd gnd cell_6t
Xbit_r105_c211 bl_211 br_211 wl_105 vdd gnd cell_6t
Xbit_r106_c211 bl_211 br_211 wl_106 vdd gnd cell_6t
Xbit_r107_c211 bl_211 br_211 wl_107 vdd gnd cell_6t
Xbit_r108_c211 bl_211 br_211 wl_108 vdd gnd cell_6t
Xbit_r109_c211 bl_211 br_211 wl_109 vdd gnd cell_6t
Xbit_r110_c211 bl_211 br_211 wl_110 vdd gnd cell_6t
Xbit_r111_c211 bl_211 br_211 wl_111 vdd gnd cell_6t
Xbit_r112_c211 bl_211 br_211 wl_112 vdd gnd cell_6t
Xbit_r113_c211 bl_211 br_211 wl_113 vdd gnd cell_6t
Xbit_r114_c211 bl_211 br_211 wl_114 vdd gnd cell_6t
Xbit_r115_c211 bl_211 br_211 wl_115 vdd gnd cell_6t
Xbit_r116_c211 bl_211 br_211 wl_116 vdd gnd cell_6t
Xbit_r117_c211 bl_211 br_211 wl_117 vdd gnd cell_6t
Xbit_r118_c211 bl_211 br_211 wl_118 vdd gnd cell_6t
Xbit_r119_c211 bl_211 br_211 wl_119 vdd gnd cell_6t
Xbit_r120_c211 bl_211 br_211 wl_120 vdd gnd cell_6t
Xbit_r121_c211 bl_211 br_211 wl_121 vdd gnd cell_6t
Xbit_r122_c211 bl_211 br_211 wl_122 vdd gnd cell_6t
Xbit_r123_c211 bl_211 br_211 wl_123 vdd gnd cell_6t
Xbit_r124_c211 bl_211 br_211 wl_124 vdd gnd cell_6t
Xbit_r125_c211 bl_211 br_211 wl_125 vdd gnd cell_6t
Xbit_r126_c211 bl_211 br_211 wl_126 vdd gnd cell_6t
Xbit_r127_c211 bl_211 br_211 wl_127 vdd gnd cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd cell_6t
Xbit_r1_c212 bl_212 br_212 wl_1 vdd gnd cell_6t
Xbit_r2_c212 bl_212 br_212 wl_2 vdd gnd cell_6t
Xbit_r3_c212 bl_212 br_212 wl_3 vdd gnd cell_6t
Xbit_r4_c212 bl_212 br_212 wl_4 vdd gnd cell_6t
Xbit_r5_c212 bl_212 br_212 wl_5 vdd gnd cell_6t
Xbit_r6_c212 bl_212 br_212 wl_6 vdd gnd cell_6t
Xbit_r7_c212 bl_212 br_212 wl_7 vdd gnd cell_6t
Xbit_r8_c212 bl_212 br_212 wl_8 vdd gnd cell_6t
Xbit_r9_c212 bl_212 br_212 wl_9 vdd gnd cell_6t
Xbit_r10_c212 bl_212 br_212 wl_10 vdd gnd cell_6t
Xbit_r11_c212 bl_212 br_212 wl_11 vdd gnd cell_6t
Xbit_r12_c212 bl_212 br_212 wl_12 vdd gnd cell_6t
Xbit_r13_c212 bl_212 br_212 wl_13 vdd gnd cell_6t
Xbit_r14_c212 bl_212 br_212 wl_14 vdd gnd cell_6t
Xbit_r15_c212 bl_212 br_212 wl_15 vdd gnd cell_6t
Xbit_r16_c212 bl_212 br_212 wl_16 vdd gnd cell_6t
Xbit_r17_c212 bl_212 br_212 wl_17 vdd gnd cell_6t
Xbit_r18_c212 bl_212 br_212 wl_18 vdd gnd cell_6t
Xbit_r19_c212 bl_212 br_212 wl_19 vdd gnd cell_6t
Xbit_r20_c212 bl_212 br_212 wl_20 vdd gnd cell_6t
Xbit_r21_c212 bl_212 br_212 wl_21 vdd gnd cell_6t
Xbit_r22_c212 bl_212 br_212 wl_22 vdd gnd cell_6t
Xbit_r23_c212 bl_212 br_212 wl_23 vdd gnd cell_6t
Xbit_r24_c212 bl_212 br_212 wl_24 vdd gnd cell_6t
Xbit_r25_c212 bl_212 br_212 wl_25 vdd gnd cell_6t
Xbit_r26_c212 bl_212 br_212 wl_26 vdd gnd cell_6t
Xbit_r27_c212 bl_212 br_212 wl_27 vdd gnd cell_6t
Xbit_r28_c212 bl_212 br_212 wl_28 vdd gnd cell_6t
Xbit_r29_c212 bl_212 br_212 wl_29 vdd gnd cell_6t
Xbit_r30_c212 bl_212 br_212 wl_30 vdd gnd cell_6t
Xbit_r31_c212 bl_212 br_212 wl_31 vdd gnd cell_6t
Xbit_r32_c212 bl_212 br_212 wl_32 vdd gnd cell_6t
Xbit_r33_c212 bl_212 br_212 wl_33 vdd gnd cell_6t
Xbit_r34_c212 bl_212 br_212 wl_34 vdd gnd cell_6t
Xbit_r35_c212 bl_212 br_212 wl_35 vdd gnd cell_6t
Xbit_r36_c212 bl_212 br_212 wl_36 vdd gnd cell_6t
Xbit_r37_c212 bl_212 br_212 wl_37 vdd gnd cell_6t
Xbit_r38_c212 bl_212 br_212 wl_38 vdd gnd cell_6t
Xbit_r39_c212 bl_212 br_212 wl_39 vdd gnd cell_6t
Xbit_r40_c212 bl_212 br_212 wl_40 vdd gnd cell_6t
Xbit_r41_c212 bl_212 br_212 wl_41 vdd gnd cell_6t
Xbit_r42_c212 bl_212 br_212 wl_42 vdd gnd cell_6t
Xbit_r43_c212 bl_212 br_212 wl_43 vdd gnd cell_6t
Xbit_r44_c212 bl_212 br_212 wl_44 vdd gnd cell_6t
Xbit_r45_c212 bl_212 br_212 wl_45 vdd gnd cell_6t
Xbit_r46_c212 bl_212 br_212 wl_46 vdd gnd cell_6t
Xbit_r47_c212 bl_212 br_212 wl_47 vdd gnd cell_6t
Xbit_r48_c212 bl_212 br_212 wl_48 vdd gnd cell_6t
Xbit_r49_c212 bl_212 br_212 wl_49 vdd gnd cell_6t
Xbit_r50_c212 bl_212 br_212 wl_50 vdd gnd cell_6t
Xbit_r51_c212 bl_212 br_212 wl_51 vdd gnd cell_6t
Xbit_r52_c212 bl_212 br_212 wl_52 vdd gnd cell_6t
Xbit_r53_c212 bl_212 br_212 wl_53 vdd gnd cell_6t
Xbit_r54_c212 bl_212 br_212 wl_54 vdd gnd cell_6t
Xbit_r55_c212 bl_212 br_212 wl_55 vdd gnd cell_6t
Xbit_r56_c212 bl_212 br_212 wl_56 vdd gnd cell_6t
Xbit_r57_c212 bl_212 br_212 wl_57 vdd gnd cell_6t
Xbit_r58_c212 bl_212 br_212 wl_58 vdd gnd cell_6t
Xbit_r59_c212 bl_212 br_212 wl_59 vdd gnd cell_6t
Xbit_r60_c212 bl_212 br_212 wl_60 vdd gnd cell_6t
Xbit_r61_c212 bl_212 br_212 wl_61 vdd gnd cell_6t
Xbit_r62_c212 bl_212 br_212 wl_62 vdd gnd cell_6t
Xbit_r63_c212 bl_212 br_212 wl_63 vdd gnd cell_6t
Xbit_r64_c212 bl_212 br_212 wl_64 vdd gnd cell_6t
Xbit_r65_c212 bl_212 br_212 wl_65 vdd gnd cell_6t
Xbit_r66_c212 bl_212 br_212 wl_66 vdd gnd cell_6t
Xbit_r67_c212 bl_212 br_212 wl_67 vdd gnd cell_6t
Xbit_r68_c212 bl_212 br_212 wl_68 vdd gnd cell_6t
Xbit_r69_c212 bl_212 br_212 wl_69 vdd gnd cell_6t
Xbit_r70_c212 bl_212 br_212 wl_70 vdd gnd cell_6t
Xbit_r71_c212 bl_212 br_212 wl_71 vdd gnd cell_6t
Xbit_r72_c212 bl_212 br_212 wl_72 vdd gnd cell_6t
Xbit_r73_c212 bl_212 br_212 wl_73 vdd gnd cell_6t
Xbit_r74_c212 bl_212 br_212 wl_74 vdd gnd cell_6t
Xbit_r75_c212 bl_212 br_212 wl_75 vdd gnd cell_6t
Xbit_r76_c212 bl_212 br_212 wl_76 vdd gnd cell_6t
Xbit_r77_c212 bl_212 br_212 wl_77 vdd gnd cell_6t
Xbit_r78_c212 bl_212 br_212 wl_78 vdd gnd cell_6t
Xbit_r79_c212 bl_212 br_212 wl_79 vdd gnd cell_6t
Xbit_r80_c212 bl_212 br_212 wl_80 vdd gnd cell_6t
Xbit_r81_c212 bl_212 br_212 wl_81 vdd gnd cell_6t
Xbit_r82_c212 bl_212 br_212 wl_82 vdd gnd cell_6t
Xbit_r83_c212 bl_212 br_212 wl_83 vdd gnd cell_6t
Xbit_r84_c212 bl_212 br_212 wl_84 vdd gnd cell_6t
Xbit_r85_c212 bl_212 br_212 wl_85 vdd gnd cell_6t
Xbit_r86_c212 bl_212 br_212 wl_86 vdd gnd cell_6t
Xbit_r87_c212 bl_212 br_212 wl_87 vdd gnd cell_6t
Xbit_r88_c212 bl_212 br_212 wl_88 vdd gnd cell_6t
Xbit_r89_c212 bl_212 br_212 wl_89 vdd gnd cell_6t
Xbit_r90_c212 bl_212 br_212 wl_90 vdd gnd cell_6t
Xbit_r91_c212 bl_212 br_212 wl_91 vdd gnd cell_6t
Xbit_r92_c212 bl_212 br_212 wl_92 vdd gnd cell_6t
Xbit_r93_c212 bl_212 br_212 wl_93 vdd gnd cell_6t
Xbit_r94_c212 bl_212 br_212 wl_94 vdd gnd cell_6t
Xbit_r95_c212 bl_212 br_212 wl_95 vdd gnd cell_6t
Xbit_r96_c212 bl_212 br_212 wl_96 vdd gnd cell_6t
Xbit_r97_c212 bl_212 br_212 wl_97 vdd gnd cell_6t
Xbit_r98_c212 bl_212 br_212 wl_98 vdd gnd cell_6t
Xbit_r99_c212 bl_212 br_212 wl_99 vdd gnd cell_6t
Xbit_r100_c212 bl_212 br_212 wl_100 vdd gnd cell_6t
Xbit_r101_c212 bl_212 br_212 wl_101 vdd gnd cell_6t
Xbit_r102_c212 bl_212 br_212 wl_102 vdd gnd cell_6t
Xbit_r103_c212 bl_212 br_212 wl_103 vdd gnd cell_6t
Xbit_r104_c212 bl_212 br_212 wl_104 vdd gnd cell_6t
Xbit_r105_c212 bl_212 br_212 wl_105 vdd gnd cell_6t
Xbit_r106_c212 bl_212 br_212 wl_106 vdd gnd cell_6t
Xbit_r107_c212 bl_212 br_212 wl_107 vdd gnd cell_6t
Xbit_r108_c212 bl_212 br_212 wl_108 vdd gnd cell_6t
Xbit_r109_c212 bl_212 br_212 wl_109 vdd gnd cell_6t
Xbit_r110_c212 bl_212 br_212 wl_110 vdd gnd cell_6t
Xbit_r111_c212 bl_212 br_212 wl_111 vdd gnd cell_6t
Xbit_r112_c212 bl_212 br_212 wl_112 vdd gnd cell_6t
Xbit_r113_c212 bl_212 br_212 wl_113 vdd gnd cell_6t
Xbit_r114_c212 bl_212 br_212 wl_114 vdd gnd cell_6t
Xbit_r115_c212 bl_212 br_212 wl_115 vdd gnd cell_6t
Xbit_r116_c212 bl_212 br_212 wl_116 vdd gnd cell_6t
Xbit_r117_c212 bl_212 br_212 wl_117 vdd gnd cell_6t
Xbit_r118_c212 bl_212 br_212 wl_118 vdd gnd cell_6t
Xbit_r119_c212 bl_212 br_212 wl_119 vdd gnd cell_6t
Xbit_r120_c212 bl_212 br_212 wl_120 vdd gnd cell_6t
Xbit_r121_c212 bl_212 br_212 wl_121 vdd gnd cell_6t
Xbit_r122_c212 bl_212 br_212 wl_122 vdd gnd cell_6t
Xbit_r123_c212 bl_212 br_212 wl_123 vdd gnd cell_6t
Xbit_r124_c212 bl_212 br_212 wl_124 vdd gnd cell_6t
Xbit_r125_c212 bl_212 br_212 wl_125 vdd gnd cell_6t
Xbit_r126_c212 bl_212 br_212 wl_126 vdd gnd cell_6t
Xbit_r127_c212 bl_212 br_212 wl_127 vdd gnd cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd cell_6t
Xbit_r1_c213 bl_213 br_213 wl_1 vdd gnd cell_6t
Xbit_r2_c213 bl_213 br_213 wl_2 vdd gnd cell_6t
Xbit_r3_c213 bl_213 br_213 wl_3 vdd gnd cell_6t
Xbit_r4_c213 bl_213 br_213 wl_4 vdd gnd cell_6t
Xbit_r5_c213 bl_213 br_213 wl_5 vdd gnd cell_6t
Xbit_r6_c213 bl_213 br_213 wl_6 vdd gnd cell_6t
Xbit_r7_c213 bl_213 br_213 wl_7 vdd gnd cell_6t
Xbit_r8_c213 bl_213 br_213 wl_8 vdd gnd cell_6t
Xbit_r9_c213 bl_213 br_213 wl_9 vdd gnd cell_6t
Xbit_r10_c213 bl_213 br_213 wl_10 vdd gnd cell_6t
Xbit_r11_c213 bl_213 br_213 wl_11 vdd gnd cell_6t
Xbit_r12_c213 bl_213 br_213 wl_12 vdd gnd cell_6t
Xbit_r13_c213 bl_213 br_213 wl_13 vdd gnd cell_6t
Xbit_r14_c213 bl_213 br_213 wl_14 vdd gnd cell_6t
Xbit_r15_c213 bl_213 br_213 wl_15 vdd gnd cell_6t
Xbit_r16_c213 bl_213 br_213 wl_16 vdd gnd cell_6t
Xbit_r17_c213 bl_213 br_213 wl_17 vdd gnd cell_6t
Xbit_r18_c213 bl_213 br_213 wl_18 vdd gnd cell_6t
Xbit_r19_c213 bl_213 br_213 wl_19 vdd gnd cell_6t
Xbit_r20_c213 bl_213 br_213 wl_20 vdd gnd cell_6t
Xbit_r21_c213 bl_213 br_213 wl_21 vdd gnd cell_6t
Xbit_r22_c213 bl_213 br_213 wl_22 vdd gnd cell_6t
Xbit_r23_c213 bl_213 br_213 wl_23 vdd gnd cell_6t
Xbit_r24_c213 bl_213 br_213 wl_24 vdd gnd cell_6t
Xbit_r25_c213 bl_213 br_213 wl_25 vdd gnd cell_6t
Xbit_r26_c213 bl_213 br_213 wl_26 vdd gnd cell_6t
Xbit_r27_c213 bl_213 br_213 wl_27 vdd gnd cell_6t
Xbit_r28_c213 bl_213 br_213 wl_28 vdd gnd cell_6t
Xbit_r29_c213 bl_213 br_213 wl_29 vdd gnd cell_6t
Xbit_r30_c213 bl_213 br_213 wl_30 vdd gnd cell_6t
Xbit_r31_c213 bl_213 br_213 wl_31 vdd gnd cell_6t
Xbit_r32_c213 bl_213 br_213 wl_32 vdd gnd cell_6t
Xbit_r33_c213 bl_213 br_213 wl_33 vdd gnd cell_6t
Xbit_r34_c213 bl_213 br_213 wl_34 vdd gnd cell_6t
Xbit_r35_c213 bl_213 br_213 wl_35 vdd gnd cell_6t
Xbit_r36_c213 bl_213 br_213 wl_36 vdd gnd cell_6t
Xbit_r37_c213 bl_213 br_213 wl_37 vdd gnd cell_6t
Xbit_r38_c213 bl_213 br_213 wl_38 vdd gnd cell_6t
Xbit_r39_c213 bl_213 br_213 wl_39 vdd gnd cell_6t
Xbit_r40_c213 bl_213 br_213 wl_40 vdd gnd cell_6t
Xbit_r41_c213 bl_213 br_213 wl_41 vdd gnd cell_6t
Xbit_r42_c213 bl_213 br_213 wl_42 vdd gnd cell_6t
Xbit_r43_c213 bl_213 br_213 wl_43 vdd gnd cell_6t
Xbit_r44_c213 bl_213 br_213 wl_44 vdd gnd cell_6t
Xbit_r45_c213 bl_213 br_213 wl_45 vdd gnd cell_6t
Xbit_r46_c213 bl_213 br_213 wl_46 vdd gnd cell_6t
Xbit_r47_c213 bl_213 br_213 wl_47 vdd gnd cell_6t
Xbit_r48_c213 bl_213 br_213 wl_48 vdd gnd cell_6t
Xbit_r49_c213 bl_213 br_213 wl_49 vdd gnd cell_6t
Xbit_r50_c213 bl_213 br_213 wl_50 vdd gnd cell_6t
Xbit_r51_c213 bl_213 br_213 wl_51 vdd gnd cell_6t
Xbit_r52_c213 bl_213 br_213 wl_52 vdd gnd cell_6t
Xbit_r53_c213 bl_213 br_213 wl_53 vdd gnd cell_6t
Xbit_r54_c213 bl_213 br_213 wl_54 vdd gnd cell_6t
Xbit_r55_c213 bl_213 br_213 wl_55 vdd gnd cell_6t
Xbit_r56_c213 bl_213 br_213 wl_56 vdd gnd cell_6t
Xbit_r57_c213 bl_213 br_213 wl_57 vdd gnd cell_6t
Xbit_r58_c213 bl_213 br_213 wl_58 vdd gnd cell_6t
Xbit_r59_c213 bl_213 br_213 wl_59 vdd gnd cell_6t
Xbit_r60_c213 bl_213 br_213 wl_60 vdd gnd cell_6t
Xbit_r61_c213 bl_213 br_213 wl_61 vdd gnd cell_6t
Xbit_r62_c213 bl_213 br_213 wl_62 vdd gnd cell_6t
Xbit_r63_c213 bl_213 br_213 wl_63 vdd gnd cell_6t
Xbit_r64_c213 bl_213 br_213 wl_64 vdd gnd cell_6t
Xbit_r65_c213 bl_213 br_213 wl_65 vdd gnd cell_6t
Xbit_r66_c213 bl_213 br_213 wl_66 vdd gnd cell_6t
Xbit_r67_c213 bl_213 br_213 wl_67 vdd gnd cell_6t
Xbit_r68_c213 bl_213 br_213 wl_68 vdd gnd cell_6t
Xbit_r69_c213 bl_213 br_213 wl_69 vdd gnd cell_6t
Xbit_r70_c213 bl_213 br_213 wl_70 vdd gnd cell_6t
Xbit_r71_c213 bl_213 br_213 wl_71 vdd gnd cell_6t
Xbit_r72_c213 bl_213 br_213 wl_72 vdd gnd cell_6t
Xbit_r73_c213 bl_213 br_213 wl_73 vdd gnd cell_6t
Xbit_r74_c213 bl_213 br_213 wl_74 vdd gnd cell_6t
Xbit_r75_c213 bl_213 br_213 wl_75 vdd gnd cell_6t
Xbit_r76_c213 bl_213 br_213 wl_76 vdd gnd cell_6t
Xbit_r77_c213 bl_213 br_213 wl_77 vdd gnd cell_6t
Xbit_r78_c213 bl_213 br_213 wl_78 vdd gnd cell_6t
Xbit_r79_c213 bl_213 br_213 wl_79 vdd gnd cell_6t
Xbit_r80_c213 bl_213 br_213 wl_80 vdd gnd cell_6t
Xbit_r81_c213 bl_213 br_213 wl_81 vdd gnd cell_6t
Xbit_r82_c213 bl_213 br_213 wl_82 vdd gnd cell_6t
Xbit_r83_c213 bl_213 br_213 wl_83 vdd gnd cell_6t
Xbit_r84_c213 bl_213 br_213 wl_84 vdd gnd cell_6t
Xbit_r85_c213 bl_213 br_213 wl_85 vdd gnd cell_6t
Xbit_r86_c213 bl_213 br_213 wl_86 vdd gnd cell_6t
Xbit_r87_c213 bl_213 br_213 wl_87 vdd gnd cell_6t
Xbit_r88_c213 bl_213 br_213 wl_88 vdd gnd cell_6t
Xbit_r89_c213 bl_213 br_213 wl_89 vdd gnd cell_6t
Xbit_r90_c213 bl_213 br_213 wl_90 vdd gnd cell_6t
Xbit_r91_c213 bl_213 br_213 wl_91 vdd gnd cell_6t
Xbit_r92_c213 bl_213 br_213 wl_92 vdd gnd cell_6t
Xbit_r93_c213 bl_213 br_213 wl_93 vdd gnd cell_6t
Xbit_r94_c213 bl_213 br_213 wl_94 vdd gnd cell_6t
Xbit_r95_c213 bl_213 br_213 wl_95 vdd gnd cell_6t
Xbit_r96_c213 bl_213 br_213 wl_96 vdd gnd cell_6t
Xbit_r97_c213 bl_213 br_213 wl_97 vdd gnd cell_6t
Xbit_r98_c213 bl_213 br_213 wl_98 vdd gnd cell_6t
Xbit_r99_c213 bl_213 br_213 wl_99 vdd gnd cell_6t
Xbit_r100_c213 bl_213 br_213 wl_100 vdd gnd cell_6t
Xbit_r101_c213 bl_213 br_213 wl_101 vdd gnd cell_6t
Xbit_r102_c213 bl_213 br_213 wl_102 vdd gnd cell_6t
Xbit_r103_c213 bl_213 br_213 wl_103 vdd gnd cell_6t
Xbit_r104_c213 bl_213 br_213 wl_104 vdd gnd cell_6t
Xbit_r105_c213 bl_213 br_213 wl_105 vdd gnd cell_6t
Xbit_r106_c213 bl_213 br_213 wl_106 vdd gnd cell_6t
Xbit_r107_c213 bl_213 br_213 wl_107 vdd gnd cell_6t
Xbit_r108_c213 bl_213 br_213 wl_108 vdd gnd cell_6t
Xbit_r109_c213 bl_213 br_213 wl_109 vdd gnd cell_6t
Xbit_r110_c213 bl_213 br_213 wl_110 vdd gnd cell_6t
Xbit_r111_c213 bl_213 br_213 wl_111 vdd gnd cell_6t
Xbit_r112_c213 bl_213 br_213 wl_112 vdd gnd cell_6t
Xbit_r113_c213 bl_213 br_213 wl_113 vdd gnd cell_6t
Xbit_r114_c213 bl_213 br_213 wl_114 vdd gnd cell_6t
Xbit_r115_c213 bl_213 br_213 wl_115 vdd gnd cell_6t
Xbit_r116_c213 bl_213 br_213 wl_116 vdd gnd cell_6t
Xbit_r117_c213 bl_213 br_213 wl_117 vdd gnd cell_6t
Xbit_r118_c213 bl_213 br_213 wl_118 vdd gnd cell_6t
Xbit_r119_c213 bl_213 br_213 wl_119 vdd gnd cell_6t
Xbit_r120_c213 bl_213 br_213 wl_120 vdd gnd cell_6t
Xbit_r121_c213 bl_213 br_213 wl_121 vdd gnd cell_6t
Xbit_r122_c213 bl_213 br_213 wl_122 vdd gnd cell_6t
Xbit_r123_c213 bl_213 br_213 wl_123 vdd gnd cell_6t
Xbit_r124_c213 bl_213 br_213 wl_124 vdd gnd cell_6t
Xbit_r125_c213 bl_213 br_213 wl_125 vdd gnd cell_6t
Xbit_r126_c213 bl_213 br_213 wl_126 vdd gnd cell_6t
Xbit_r127_c213 bl_213 br_213 wl_127 vdd gnd cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd cell_6t
Xbit_r1_c214 bl_214 br_214 wl_1 vdd gnd cell_6t
Xbit_r2_c214 bl_214 br_214 wl_2 vdd gnd cell_6t
Xbit_r3_c214 bl_214 br_214 wl_3 vdd gnd cell_6t
Xbit_r4_c214 bl_214 br_214 wl_4 vdd gnd cell_6t
Xbit_r5_c214 bl_214 br_214 wl_5 vdd gnd cell_6t
Xbit_r6_c214 bl_214 br_214 wl_6 vdd gnd cell_6t
Xbit_r7_c214 bl_214 br_214 wl_7 vdd gnd cell_6t
Xbit_r8_c214 bl_214 br_214 wl_8 vdd gnd cell_6t
Xbit_r9_c214 bl_214 br_214 wl_9 vdd gnd cell_6t
Xbit_r10_c214 bl_214 br_214 wl_10 vdd gnd cell_6t
Xbit_r11_c214 bl_214 br_214 wl_11 vdd gnd cell_6t
Xbit_r12_c214 bl_214 br_214 wl_12 vdd gnd cell_6t
Xbit_r13_c214 bl_214 br_214 wl_13 vdd gnd cell_6t
Xbit_r14_c214 bl_214 br_214 wl_14 vdd gnd cell_6t
Xbit_r15_c214 bl_214 br_214 wl_15 vdd gnd cell_6t
Xbit_r16_c214 bl_214 br_214 wl_16 vdd gnd cell_6t
Xbit_r17_c214 bl_214 br_214 wl_17 vdd gnd cell_6t
Xbit_r18_c214 bl_214 br_214 wl_18 vdd gnd cell_6t
Xbit_r19_c214 bl_214 br_214 wl_19 vdd gnd cell_6t
Xbit_r20_c214 bl_214 br_214 wl_20 vdd gnd cell_6t
Xbit_r21_c214 bl_214 br_214 wl_21 vdd gnd cell_6t
Xbit_r22_c214 bl_214 br_214 wl_22 vdd gnd cell_6t
Xbit_r23_c214 bl_214 br_214 wl_23 vdd gnd cell_6t
Xbit_r24_c214 bl_214 br_214 wl_24 vdd gnd cell_6t
Xbit_r25_c214 bl_214 br_214 wl_25 vdd gnd cell_6t
Xbit_r26_c214 bl_214 br_214 wl_26 vdd gnd cell_6t
Xbit_r27_c214 bl_214 br_214 wl_27 vdd gnd cell_6t
Xbit_r28_c214 bl_214 br_214 wl_28 vdd gnd cell_6t
Xbit_r29_c214 bl_214 br_214 wl_29 vdd gnd cell_6t
Xbit_r30_c214 bl_214 br_214 wl_30 vdd gnd cell_6t
Xbit_r31_c214 bl_214 br_214 wl_31 vdd gnd cell_6t
Xbit_r32_c214 bl_214 br_214 wl_32 vdd gnd cell_6t
Xbit_r33_c214 bl_214 br_214 wl_33 vdd gnd cell_6t
Xbit_r34_c214 bl_214 br_214 wl_34 vdd gnd cell_6t
Xbit_r35_c214 bl_214 br_214 wl_35 vdd gnd cell_6t
Xbit_r36_c214 bl_214 br_214 wl_36 vdd gnd cell_6t
Xbit_r37_c214 bl_214 br_214 wl_37 vdd gnd cell_6t
Xbit_r38_c214 bl_214 br_214 wl_38 vdd gnd cell_6t
Xbit_r39_c214 bl_214 br_214 wl_39 vdd gnd cell_6t
Xbit_r40_c214 bl_214 br_214 wl_40 vdd gnd cell_6t
Xbit_r41_c214 bl_214 br_214 wl_41 vdd gnd cell_6t
Xbit_r42_c214 bl_214 br_214 wl_42 vdd gnd cell_6t
Xbit_r43_c214 bl_214 br_214 wl_43 vdd gnd cell_6t
Xbit_r44_c214 bl_214 br_214 wl_44 vdd gnd cell_6t
Xbit_r45_c214 bl_214 br_214 wl_45 vdd gnd cell_6t
Xbit_r46_c214 bl_214 br_214 wl_46 vdd gnd cell_6t
Xbit_r47_c214 bl_214 br_214 wl_47 vdd gnd cell_6t
Xbit_r48_c214 bl_214 br_214 wl_48 vdd gnd cell_6t
Xbit_r49_c214 bl_214 br_214 wl_49 vdd gnd cell_6t
Xbit_r50_c214 bl_214 br_214 wl_50 vdd gnd cell_6t
Xbit_r51_c214 bl_214 br_214 wl_51 vdd gnd cell_6t
Xbit_r52_c214 bl_214 br_214 wl_52 vdd gnd cell_6t
Xbit_r53_c214 bl_214 br_214 wl_53 vdd gnd cell_6t
Xbit_r54_c214 bl_214 br_214 wl_54 vdd gnd cell_6t
Xbit_r55_c214 bl_214 br_214 wl_55 vdd gnd cell_6t
Xbit_r56_c214 bl_214 br_214 wl_56 vdd gnd cell_6t
Xbit_r57_c214 bl_214 br_214 wl_57 vdd gnd cell_6t
Xbit_r58_c214 bl_214 br_214 wl_58 vdd gnd cell_6t
Xbit_r59_c214 bl_214 br_214 wl_59 vdd gnd cell_6t
Xbit_r60_c214 bl_214 br_214 wl_60 vdd gnd cell_6t
Xbit_r61_c214 bl_214 br_214 wl_61 vdd gnd cell_6t
Xbit_r62_c214 bl_214 br_214 wl_62 vdd gnd cell_6t
Xbit_r63_c214 bl_214 br_214 wl_63 vdd gnd cell_6t
Xbit_r64_c214 bl_214 br_214 wl_64 vdd gnd cell_6t
Xbit_r65_c214 bl_214 br_214 wl_65 vdd gnd cell_6t
Xbit_r66_c214 bl_214 br_214 wl_66 vdd gnd cell_6t
Xbit_r67_c214 bl_214 br_214 wl_67 vdd gnd cell_6t
Xbit_r68_c214 bl_214 br_214 wl_68 vdd gnd cell_6t
Xbit_r69_c214 bl_214 br_214 wl_69 vdd gnd cell_6t
Xbit_r70_c214 bl_214 br_214 wl_70 vdd gnd cell_6t
Xbit_r71_c214 bl_214 br_214 wl_71 vdd gnd cell_6t
Xbit_r72_c214 bl_214 br_214 wl_72 vdd gnd cell_6t
Xbit_r73_c214 bl_214 br_214 wl_73 vdd gnd cell_6t
Xbit_r74_c214 bl_214 br_214 wl_74 vdd gnd cell_6t
Xbit_r75_c214 bl_214 br_214 wl_75 vdd gnd cell_6t
Xbit_r76_c214 bl_214 br_214 wl_76 vdd gnd cell_6t
Xbit_r77_c214 bl_214 br_214 wl_77 vdd gnd cell_6t
Xbit_r78_c214 bl_214 br_214 wl_78 vdd gnd cell_6t
Xbit_r79_c214 bl_214 br_214 wl_79 vdd gnd cell_6t
Xbit_r80_c214 bl_214 br_214 wl_80 vdd gnd cell_6t
Xbit_r81_c214 bl_214 br_214 wl_81 vdd gnd cell_6t
Xbit_r82_c214 bl_214 br_214 wl_82 vdd gnd cell_6t
Xbit_r83_c214 bl_214 br_214 wl_83 vdd gnd cell_6t
Xbit_r84_c214 bl_214 br_214 wl_84 vdd gnd cell_6t
Xbit_r85_c214 bl_214 br_214 wl_85 vdd gnd cell_6t
Xbit_r86_c214 bl_214 br_214 wl_86 vdd gnd cell_6t
Xbit_r87_c214 bl_214 br_214 wl_87 vdd gnd cell_6t
Xbit_r88_c214 bl_214 br_214 wl_88 vdd gnd cell_6t
Xbit_r89_c214 bl_214 br_214 wl_89 vdd gnd cell_6t
Xbit_r90_c214 bl_214 br_214 wl_90 vdd gnd cell_6t
Xbit_r91_c214 bl_214 br_214 wl_91 vdd gnd cell_6t
Xbit_r92_c214 bl_214 br_214 wl_92 vdd gnd cell_6t
Xbit_r93_c214 bl_214 br_214 wl_93 vdd gnd cell_6t
Xbit_r94_c214 bl_214 br_214 wl_94 vdd gnd cell_6t
Xbit_r95_c214 bl_214 br_214 wl_95 vdd gnd cell_6t
Xbit_r96_c214 bl_214 br_214 wl_96 vdd gnd cell_6t
Xbit_r97_c214 bl_214 br_214 wl_97 vdd gnd cell_6t
Xbit_r98_c214 bl_214 br_214 wl_98 vdd gnd cell_6t
Xbit_r99_c214 bl_214 br_214 wl_99 vdd gnd cell_6t
Xbit_r100_c214 bl_214 br_214 wl_100 vdd gnd cell_6t
Xbit_r101_c214 bl_214 br_214 wl_101 vdd gnd cell_6t
Xbit_r102_c214 bl_214 br_214 wl_102 vdd gnd cell_6t
Xbit_r103_c214 bl_214 br_214 wl_103 vdd gnd cell_6t
Xbit_r104_c214 bl_214 br_214 wl_104 vdd gnd cell_6t
Xbit_r105_c214 bl_214 br_214 wl_105 vdd gnd cell_6t
Xbit_r106_c214 bl_214 br_214 wl_106 vdd gnd cell_6t
Xbit_r107_c214 bl_214 br_214 wl_107 vdd gnd cell_6t
Xbit_r108_c214 bl_214 br_214 wl_108 vdd gnd cell_6t
Xbit_r109_c214 bl_214 br_214 wl_109 vdd gnd cell_6t
Xbit_r110_c214 bl_214 br_214 wl_110 vdd gnd cell_6t
Xbit_r111_c214 bl_214 br_214 wl_111 vdd gnd cell_6t
Xbit_r112_c214 bl_214 br_214 wl_112 vdd gnd cell_6t
Xbit_r113_c214 bl_214 br_214 wl_113 vdd gnd cell_6t
Xbit_r114_c214 bl_214 br_214 wl_114 vdd gnd cell_6t
Xbit_r115_c214 bl_214 br_214 wl_115 vdd gnd cell_6t
Xbit_r116_c214 bl_214 br_214 wl_116 vdd gnd cell_6t
Xbit_r117_c214 bl_214 br_214 wl_117 vdd gnd cell_6t
Xbit_r118_c214 bl_214 br_214 wl_118 vdd gnd cell_6t
Xbit_r119_c214 bl_214 br_214 wl_119 vdd gnd cell_6t
Xbit_r120_c214 bl_214 br_214 wl_120 vdd gnd cell_6t
Xbit_r121_c214 bl_214 br_214 wl_121 vdd gnd cell_6t
Xbit_r122_c214 bl_214 br_214 wl_122 vdd gnd cell_6t
Xbit_r123_c214 bl_214 br_214 wl_123 vdd gnd cell_6t
Xbit_r124_c214 bl_214 br_214 wl_124 vdd gnd cell_6t
Xbit_r125_c214 bl_214 br_214 wl_125 vdd gnd cell_6t
Xbit_r126_c214 bl_214 br_214 wl_126 vdd gnd cell_6t
Xbit_r127_c214 bl_214 br_214 wl_127 vdd gnd cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd cell_6t
Xbit_r1_c215 bl_215 br_215 wl_1 vdd gnd cell_6t
Xbit_r2_c215 bl_215 br_215 wl_2 vdd gnd cell_6t
Xbit_r3_c215 bl_215 br_215 wl_3 vdd gnd cell_6t
Xbit_r4_c215 bl_215 br_215 wl_4 vdd gnd cell_6t
Xbit_r5_c215 bl_215 br_215 wl_5 vdd gnd cell_6t
Xbit_r6_c215 bl_215 br_215 wl_6 vdd gnd cell_6t
Xbit_r7_c215 bl_215 br_215 wl_7 vdd gnd cell_6t
Xbit_r8_c215 bl_215 br_215 wl_8 vdd gnd cell_6t
Xbit_r9_c215 bl_215 br_215 wl_9 vdd gnd cell_6t
Xbit_r10_c215 bl_215 br_215 wl_10 vdd gnd cell_6t
Xbit_r11_c215 bl_215 br_215 wl_11 vdd gnd cell_6t
Xbit_r12_c215 bl_215 br_215 wl_12 vdd gnd cell_6t
Xbit_r13_c215 bl_215 br_215 wl_13 vdd gnd cell_6t
Xbit_r14_c215 bl_215 br_215 wl_14 vdd gnd cell_6t
Xbit_r15_c215 bl_215 br_215 wl_15 vdd gnd cell_6t
Xbit_r16_c215 bl_215 br_215 wl_16 vdd gnd cell_6t
Xbit_r17_c215 bl_215 br_215 wl_17 vdd gnd cell_6t
Xbit_r18_c215 bl_215 br_215 wl_18 vdd gnd cell_6t
Xbit_r19_c215 bl_215 br_215 wl_19 vdd gnd cell_6t
Xbit_r20_c215 bl_215 br_215 wl_20 vdd gnd cell_6t
Xbit_r21_c215 bl_215 br_215 wl_21 vdd gnd cell_6t
Xbit_r22_c215 bl_215 br_215 wl_22 vdd gnd cell_6t
Xbit_r23_c215 bl_215 br_215 wl_23 vdd gnd cell_6t
Xbit_r24_c215 bl_215 br_215 wl_24 vdd gnd cell_6t
Xbit_r25_c215 bl_215 br_215 wl_25 vdd gnd cell_6t
Xbit_r26_c215 bl_215 br_215 wl_26 vdd gnd cell_6t
Xbit_r27_c215 bl_215 br_215 wl_27 vdd gnd cell_6t
Xbit_r28_c215 bl_215 br_215 wl_28 vdd gnd cell_6t
Xbit_r29_c215 bl_215 br_215 wl_29 vdd gnd cell_6t
Xbit_r30_c215 bl_215 br_215 wl_30 vdd gnd cell_6t
Xbit_r31_c215 bl_215 br_215 wl_31 vdd gnd cell_6t
Xbit_r32_c215 bl_215 br_215 wl_32 vdd gnd cell_6t
Xbit_r33_c215 bl_215 br_215 wl_33 vdd gnd cell_6t
Xbit_r34_c215 bl_215 br_215 wl_34 vdd gnd cell_6t
Xbit_r35_c215 bl_215 br_215 wl_35 vdd gnd cell_6t
Xbit_r36_c215 bl_215 br_215 wl_36 vdd gnd cell_6t
Xbit_r37_c215 bl_215 br_215 wl_37 vdd gnd cell_6t
Xbit_r38_c215 bl_215 br_215 wl_38 vdd gnd cell_6t
Xbit_r39_c215 bl_215 br_215 wl_39 vdd gnd cell_6t
Xbit_r40_c215 bl_215 br_215 wl_40 vdd gnd cell_6t
Xbit_r41_c215 bl_215 br_215 wl_41 vdd gnd cell_6t
Xbit_r42_c215 bl_215 br_215 wl_42 vdd gnd cell_6t
Xbit_r43_c215 bl_215 br_215 wl_43 vdd gnd cell_6t
Xbit_r44_c215 bl_215 br_215 wl_44 vdd gnd cell_6t
Xbit_r45_c215 bl_215 br_215 wl_45 vdd gnd cell_6t
Xbit_r46_c215 bl_215 br_215 wl_46 vdd gnd cell_6t
Xbit_r47_c215 bl_215 br_215 wl_47 vdd gnd cell_6t
Xbit_r48_c215 bl_215 br_215 wl_48 vdd gnd cell_6t
Xbit_r49_c215 bl_215 br_215 wl_49 vdd gnd cell_6t
Xbit_r50_c215 bl_215 br_215 wl_50 vdd gnd cell_6t
Xbit_r51_c215 bl_215 br_215 wl_51 vdd gnd cell_6t
Xbit_r52_c215 bl_215 br_215 wl_52 vdd gnd cell_6t
Xbit_r53_c215 bl_215 br_215 wl_53 vdd gnd cell_6t
Xbit_r54_c215 bl_215 br_215 wl_54 vdd gnd cell_6t
Xbit_r55_c215 bl_215 br_215 wl_55 vdd gnd cell_6t
Xbit_r56_c215 bl_215 br_215 wl_56 vdd gnd cell_6t
Xbit_r57_c215 bl_215 br_215 wl_57 vdd gnd cell_6t
Xbit_r58_c215 bl_215 br_215 wl_58 vdd gnd cell_6t
Xbit_r59_c215 bl_215 br_215 wl_59 vdd gnd cell_6t
Xbit_r60_c215 bl_215 br_215 wl_60 vdd gnd cell_6t
Xbit_r61_c215 bl_215 br_215 wl_61 vdd gnd cell_6t
Xbit_r62_c215 bl_215 br_215 wl_62 vdd gnd cell_6t
Xbit_r63_c215 bl_215 br_215 wl_63 vdd gnd cell_6t
Xbit_r64_c215 bl_215 br_215 wl_64 vdd gnd cell_6t
Xbit_r65_c215 bl_215 br_215 wl_65 vdd gnd cell_6t
Xbit_r66_c215 bl_215 br_215 wl_66 vdd gnd cell_6t
Xbit_r67_c215 bl_215 br_215 wl_67 vdd gnd cell_6t
Xbit_r68_c215 bl_215 br_215 wl_68 vdd gnd cell_6t
Xbit_r69_c215 bl_215 br_215 wl_69 vdd gnd cell_6t
Xbit_r70_c215 bl_215 br_215 wl_70 vdd gnd cell_6t
Xbit_r71_c215 bl_215 br_215 wl_71 vdd gnd cell_6t
Xbit_r72_c215 bl_215 br_215 wl_72 vdd gnd cell_6t
Xbit_r73_c215 bl_215 br_215 wl_73 vdd gnd cell_6t
Xbit_r74_c215 bl_215 br_215 wl_74 vdd gnd cell_6t
Xbit_r75_c215 bl_215 br_215 wl_75 vdd gnd cell_6t
Xbit_r76_c215 bl_215 br_215 wl_76 vdd gnd cell_6t
Xbit_r77_c215 bl_215 br_215 wl_77 vdd gnd cell_6t
Xbit_r78_c215 bl_215 br_215 wl_78 vdd gnd cell_6t
Xbit_r79_c215 bl_215 br_215 wl_79 vdd gnd cell_6t
Xbit_r80_c215 bl_215 br_215 wl_80 vdd gnd cell_6t
Xbit_r81_c215 bl_215 br_215 wl_81 vdd gnd cell_6t
Xbit_r82_c215 bl_215 br_215 wl_82 vdd gnd cell_6t
Xbit_r83_c215 bl_215 br_215 wl_83 vdd gnd cell_6t
Xbit_r84_c215 bl_215 br_215 wl_84 vdd gnd cell_6t
Xbit_r85_c215 bl_215 br_215 wl_85 vdd gnd cell_6t
Xbit_r86_c215 bl_215 br_215 wl_86 vdd gnd cell_6t
Xbit_r87_c215 bl_215 br_215 wl_87 vdd gnd cell_6t
Xbit_r88_c215 bl_215 br_215 wl_88 vdd gnd cell_6t
Xbit_r89_c215 bl_215 br_215 wl_89 vdd gnd cell_6t
Xbit_r90_c215 bl_215 br_215 wl_90 vdd gnd cell_6t
Xbit_r91_c215 bl_215 br_215 wl_91 vdd gnd cell_6t
Xbit_r92_c215 bl_215 br_215 wl_92 vdd gnd cell_6t
Xbit_r93_c215 bl_215 br_215 wl_93 vdd gnd cell_6t
Xbit_r94_c215 bl_215 br_215 wl_94 vdd gnd cell_6t
Xbit_r95_c215 bl_215 br_215 wl_95 vdd gnd cell_6t
Xbit_r96_c215 bl_215 br_215 wl_96 vdd gnd cell_6t
Xbit_r97_c215 bl_215 br_215 wl_97 vdd gnd cell_6t
Xbit_r98_c215 bl_215 br_215 wl_98 vdd gnd cell_6t
Xbit_r99_c215 bl_215 br_215 wl_99 vdd gnd cell_6t
Xbit_r100_c215 bl_215 br_215 wl_100 vdd gnd cell_6t
Xbit_r101_c215 bl_215 br_215 wl_101 vdd gnd cell_6t
Xbit_r102_c215 bl_215 br_215 wl_102 vdd gnd cell_6t
Xbit_r103_c215 bl_215 br_215 wl_103 vdd gnd cell_6t
Xbit_r104_c215 bl_215 br_215 wl_104 vdd gnd cell_6t
Xbit_r105_c215 bl_215 br_215 wl_105 vdd gnd cell_6t
Xbit_r106_c215 bl_215 br_215 wl_106 vdd gnd cell_6t
Xbit_r107_c215 bl_215 br_215 wl_107 vdd gnd cell_6t
Xbit_r108_c215 bl_215 br_215 wl_108 vdd gnd cell_6t
Xbit_r109_c215 bl_215 br_215 wl_109 vdd gnd cell_6t
Xbit_r110_c215 bl_215 br_215 wl_110 vdd gnd cell_6t
Xbit_r111_c215 bl_215 br_215 wl_111 vdd gnd cell_6t
Xbit_r112_c215 bl_215 br_215 wl_112 vdd gnd cell_6t
Xbit_r113_c215 bl_215 br_215 wl_113 vdd gnd cell_6t
Xbit_r114_c215 bl_215 br_215 wl_114 vdd gnd cell_6t
Xbit_r115_c215 bl_215 br_215 wl_115 vdd gnd cell_6t
Xbit_r116_c215 bl_215 br_215 wl_116 vdd gnd cell_6t
Xbit_r117_c215 bl_215 br_215 wl_117 vdd gnd cell_6t
Xbit_r118_c215 bl_215 br_215 wl_118 vdd gnd cell_6t
Xbit_r119_c215 bl_215 br_215 wl_119 vdd gnd cell_6t
Xbit_r120_c215 bl_215 br_215 wl_120 vdd gnd cell_6t
Xbit_r121_c215 bl_215 br_215 wl_121 vdd gnd cell_6t
Xbit_r122_c215 bl_215 br_215 wl_122 vdd gnd cell_6t
Xbit_r123_c215 bl_215 br_215 wl_123 vdd gnd cell_6t
Xbit_r124_c215 bl_215 br_215 wl_124 vdd gnd cell_6t
Xbit_r125_c215 bl_215 br_215 wl_125 vdd gnd cell_6t
Xbit_r126_c215 bl_215 br_215 wl_126 vdd gnd cell_6t
Xbit_r127_c215 bl_215 br_215 wl_127 vdd gnd cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd cell_6t
Xbit_r1_c216 bl_216 br_216 wl_1 vdd gnd cell_6t
Xbit_r2_c216 bl_216 br_216 wl_2 vdd gnd cell_6t
Xbit_r3_c216 bl_216 br_216 wl_3 vdd gnd cell_6t
Xbit_r4_c216 bl_216 br_216 wl_4 vdd gnd cell_6t
Xbit_r5_c216 bl_216 br_216 wl_5 vdd gnd cell_6t
Xbit_r6_c216 bl_216 br_216 wl_6 vdd gnd cell_6t
Xbit_r7_c216 bl_216 br_216 wl_7 vdd gnd cell_6t
Xbit_r8_c216 bl_216 br_216 wl_8 vdd gnd cell_6t
Xbit_r9_c216 bl_216 br_216 wl_9 vdd gnd cell_6t
Xbit_r10_c216 bl_216 br_216 wl_10 vdd gnd cell_6t
Xbit_r11_c216 bl_216 br_216 wl_11 vdd gnd cell_6t
Xbit_r12_c216 bl_216 br_216 wl_12 vdd gnd cell_6t
Xbit_r13_c216 bl_216 br_216 wl_13 vdd gnd cell_6t
Xbit_r14_c216 bl_216 br_216 wl_14 vdd gnd cell_6t
Xbit_r15_c216 bl_216 br_216 wl_15 vdd gnd cell_6t
Xbit_r16_c216 bl_216 br_216 wl_16 vdd gnd cell_6t
Xbit_r17_c216 bl_216 br_216 wl_17 vdd gnd cell_6t
Xbit_r18_c216 bl_216 br_216 wl_18 vdd gnd cell_6t
Xbit_r19_c216 bl_216 br_216 wl_19 vdd gnd cell_6t
Xbit_r20_c216 bl_216 br_216 wl_20 vdd gnd cell_6t
Xbit_r21_c216 bl_216 br_216 wl_21 vdd gnd cell_6t
Xbit_r22_c216 bl_216 br_216 wl_22 vdd gnd cell_6t
Xbit_r23_c216 bl_216 br_216 wl_23 vdd gnd cell_6t
Xbit_r24_c216 bl_216 br_216 wl_24 vdd gnd cell_6t
Xbit_r25_c216 bl_216 br_216 wl_25 vdd gnd cell_6t
Xbit_r26_c216 bl_216 br_216 wl_26 vdd gnd cell_6t
Xbit_r27_c216 bl_216 br_216 wl_27 vdd gnd cell_6t
Xbit_r28_c216 bl_216 br_216 wl_28 vdd gnd cell_6t
Xbit_r29_c216 bl_216 br_216 wl_29 vdd gnd cell_6t
Xbit_r30_c216 bl_216 br_216 wl_30 vdd gnd cell_6t
Xbit_r31_c216 bl_216 br_216 wl_31 vdd gnd cell_6t
Xbit_r32_c216 bl_216 br_216 wl_32 vdd gnd cell_6t
Xbit_r33_c216 bl_216 br_216 wl_33 vdd gnd cell_6t
Xbit_r34_c216 bl_216 br_216 wl_34 vdd gnd cell_6t
Xbit_r35_c216 bl_216 br_216 wl_35 vdd gnd cell_6t
Xbit_r36_c216 bl_216 br_216 wl_36 vdd gnd cell_6t
Xbit_r37_c216 bl_216 br_216 wl_37 vdd gnd cell_6t
Xbit_r38_c216 bl_216 br_216 wl_38 vdd gnd cell_6t
Xbit_r39_c216 bl_216 br_216 wl_39 vdd gnd cell_6t
Xbit_r40_c216 bl_216 br_216 wl_40 vdd gnd cell_6t
Xbit_r41_c216 bl_216 br_216 wl_41 vdd gnd cell_6t
Xbit_r42_c216 bl_216 br_216 wl_42 vdd gnd cell_6t
Xbit_r43_c216 bl_216 br_216 wl_43 vdd gnd cell_6t
Xbit_r44_c216 bl_216 br_216 wl_44 vdd gnd cell_6t
Xbit_r45_c216 bl_216 br_216 wl_45 vdd gnd cell_6t
Xbit_r46_c216 bl_216 br_216 wl_46 vdd gnd cell_6t
Xbit_r47_c216 bl_216 br_216 wl_47 vdd gnd cell_6t
Xbit_r48_c216 bl_216 br_216 wl_48 vdd gnd cell_6t
Xbit_r49_c216 bl_216 br_216 wl_49 vdd gnd cell_6t
Xbit_r50_c216 bl_216 br_216 wl_50 vdd gnd cell_6t
Xbit_r51_c216 bl_216 br_216 wl_51 vdd gnd cell_6t
Xbit_r52_c216 bl_216 br_216 wl_52 vdd gnd cell_6t
Xbit_r53_c216 bl_216 br_216 wl_53 vdd gnd cell_6t
Xbit_r54_c216 bl_216 br_216 wl_54 vdd gnd cell_6t
Xbit_r55_c216 bl_216 br_216 wl_55 vdd gnd cell_6t
Xbit_r56_c216 bl_216 br_216 wl_56 vdd gnd cell_6t
Xbit_r57_c216 bl_216 br_216 wl_57 vdd gnd cell_6t
Xbit_r58_c216 bl_216 br_216 wl_58 vdd gnd cell_6t
Xbit_r59_c216 bl_216 br_216 wl_59 vdd gnd cell_6t
Xbit_r60_c216 bl_216 br_216 wl_60 vdd gnd cell_6t
Xbit_r61_c216 bl_216 br_216 wl_61 vdd gnd cell_6t
Xbit_r62_c216 bl_216 br_216 wl_62 vdd gnd cell_6t
Xbit_r63_c216 bl_216 br_216 wl_63 vdd gnd cell_6t
Xbit_r64_c216 bl_216 br_216 wl_64 vdd gnd cell_6t
Xbit_r65_c216 bl_216 br_216 wl_65 vdd gnd cell_6t
Xbit_r66_c216 bl_216 br_216 wl_66 vdd gnd cell_6t
Xbit_r67_c216 bl_216 br_216 wl_67 vdd gnd cell_6t
Xbit_r68_c216 bl_216 br_216 wl_68 vdd gnd cell_6t
Xbit_r69_c216 bl_216 br_216 wl_69 vdd gnd cell_6t
Xbit_r70_c216 bl_216 br_216 wl_70 vdd gnd cell_6t
Xbit_r71_c216 bl_216 br_216 wl_71 vdd gnd cell_6t
Xbit_r72_c216 bl_216 br_216 wl_72 vdd gnd cell_6t
Xbit_r73_c216 bl_216 br_216 wl_73 vdd gnd cell_6t
Xbit_r74_c216 bl_216 br_216 wl_74 vdd gnd cell_6t
Xbit_r75_c216 bl_216 br_216 wl_75 vdd gnd cell_6t
Xbit_r76_c216 bl_216 br_216 wl_76 vdd gnd cell_6t
Xbit_r77_c216 bl_216 br_216 wl_77 vdd gnd cell_6t
Xbit_r78_c216 bl_216 br_216 wl_78 vdd gnd cell_6t
Xbit_r79_c216 bl_216 br_216 wl_79 vdd gnd cell_6t
Xbit_r80_c216 bl_216 br_216 wl_80 vdd gnd cell_6t
Xbit_r81_c216 bl_216 br_216 wl_81 vdd gnd cell_6t
Xbit_r82_c216 bl_216 br_216 wl_82 vdd gnd cell_6t
Xbit_r83_c216 bl_216 br_216 wl_83 vdd gnd cell_6t
Xbit_r84_c216 bl_216 br_216 wl_84 vdd gnd cell_6t
Xbit_r85_c216 bl_216 br_216 wl_85 vdd gnd cell_6t
Xbit_r86_c216 bl_216 br_216 wl_86 vdd gnd cell_6t
Xbit_r87_c216 bl_216 br_216 wl_87 vdd gnd cell_6t
Xbit_r88_c216 bl_216 br_216 wl_88 vdd gnd cell_6t
Xbit_r89_c216 bl_216 br_216 wl_89 vdd gnd cell_6t
Xbit_r90_c216 bl_216 br_216 wl_90 vdd gnd cell_6t
Xbit_r91_c216 bl_216 br_216 wl_91 vdd gnd cell_6t
Xbit_r92_c216 bl_216 br_216 wl_92 vdd gnd cell_6t
Xbit_r93_c216 bl_216 br_216 wl_93 vdd gnd cell_6t
Xbit_r94_c216 bl_216 br_216 wl_94 vdd gnd cell_6t
Xbit_r95_c216 bl_216 br_216 wl_95 vdd gnd cell_6t
Xbit_r96_c216 bl_216 br_216 wl_96 vdd gnd cell_6t
Xbit_r97_c216 bl_216 br_216 wl_97 vdd gnd cell_6t
Xbit_r98_c216 bl_216 br_216 wl_98 vdd gnd cell_6t
Xbit_r99_c216 bl_216 br_216 wl_99 vdd gnd cell_6t
Xbit_r100_c216 bl_216 br_216 wl_100 vdd gnd cell_6t
Xbit_r101_c216 bl_216 br_216 wl_101 vdd gnd cell_6t
Xbit_r102_c216 bl_216 br_216 wl_102 vdd gnd cell_6t
Xbit_r103_c216 bl_216 br_216 wl_103 vdd gnd cell_6t
Xbit_r104_c216 bl_216 br_216 wl_104 vdd gnd cell_6t
Xbit_r105_c216 bl_216 br_216 wl_105 vdd gnd cell_6t
Xbit_r106_c216 bl_216 br_216 wl_106 vdd gnd cell_6t
Xbit_r107_c216 bl_216 br_216 wl_107 vdd gnd cell_6t
Xbit_r108_c216 bl_216 br_216 wl_108 vdd gnd cell_6t
Xbit_r109_c216 bl_216 br_216 wl_109 vdd gnd cell_6t
Xbit_r110_c216 bl_216 br_216 wl_110 vdd gnd cell_6t
Xbit_r111_c216 bl_216 br_216 wl_111 vdd gnd cell_6t
Xbit_r112_c216 bl_216 br_216 wl_112 vdd gnd cell_6t
Xbit_r113_c216 bl_216 br_216 wl_113 vdd gnd cell_6t
Xbit_r114_c216 bl_216 br_216 wl_114 vdd gnd cell_6t
Xbit_r115_c216 bl_216 br_216 wl_115 vdd gnd cell_6t
Xbit_r116_c216 bl_216 br_216 wl_116 vdd gnd cell_6t
Xbit_r117_c216 bl_216 br_216 wl_117 vdd gnd cell_6t
Xbit_r118_c216 bl_216 br_216 wl_118 vdd gnd cell_6t
Xbit_r119_c216 bl_216 br_216 wl_119 vdd gnd cell_6t
Xbit_r120_c216 bl_216 br_216 wl_120 vdd gnd cell_6t
Xbit_r121_c216 bl_216 br_216 wl_121 vdd gnd cell_6t
Xbit_r122_c216 bl_216 br_216 wl_122 vdd gnd cell_6t
Xbit_r123_c216 bl_216 br_216 wl_123 vdd gnd cell_6t
Xbit_r124_c216 bl_216 br_216 wl_124 vdd gnd cell_6t
Xbit_r125_c216 bl_216 br_216 wl_125 vdd gnd cell_6t
Xbit_r126_c216 bl_216 br_216 wl_126 vdd gnd cell_6t
Xbit_r127_c216 bl_216 br_216 wl_127 vdd gnd cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd cell_6t
Xbit_r1_c217 bl_217 br_217 wl_1 vdd gnd cell_6t
Xbit_r2_c217 bl_217 br_217 wl_2 vdd gnd cell_6t
Xbit_r3_c217 bl_217 br_217 wl_3 vdd gnd cell_6t
Xbit_r4_c217 bl_217 br_217 wl_4 vdd gnd cell_6t
Xbit_r5_c217 bl_217 br_217 wl_5 vdd gnd cell_6t
Xbit_r6_c217 bl_217 br_217 wl_6 vdd gnd cell_6t
Xbit_r7_c217 bl_217 br_217 wl_7 vdd gnd cell_6t
Xbit_r8_c217 bl_217 br_217 wl_8 vdd gnd cell_6t
Xbit_r9_c217 bl_217 br_217 wl_9 vdd gnd cell_6t
Xbit_r10_c217 bl_217 br_217 wl_10 vdd gnd cell_6t
Xbit_r11_c217 bl_217 br_217 wl_11 vdd gnd cell_6t
Xbit_r12_c217 bl_217 br_217 wl_12 vdd gnd cell_6t
Xbit_r13_c217 bl_217 br_217 wl_13 vdd gnd cell_6t
Xbit_r14_c217 bl_217 br_217 wl_14 vdd gnd cell_6t
Xbit_r15_c217 bl_217 br_217 wl_15 vdd gnd cell_6t
Xbit_r16_c217 bl_217 br_217 wl_16 vdd gnd cell_6t
Xbit_r17_c217 bl_217 br_217 wl_17 vdd gnd cell_6t
Xbit_r18_c217 bl_217 br_217 wl_18 vdd gnd cell_6t
Xbit_r19_c217 bl_217 br_217 wl_19 vdd gnd cell_6t
Xbit_r20_c217 bl_217 br_217 wl_20 vdd gnd cell_6t
Xbit_r21_c217 bl_217 br_217 wl_21 vdd gnd cell_6t
Xbit_r22_c217 bl_217 br_217 wl_22 vdd gnd cell_6t
Xbit_r23_c217 bl_217 br_217 wl_23 vdd gnd cell_6t
Xbit_r24_c217 bl_217 br_217 wl_24 vdd gnd cell_6t
Xbit_r25_c217 bl_217 br_217 wl_25 vdd gnd cell_6t
Xbit_r26_c217 bl_217 br_217 wl_26 vdd gnd cell_6t
Xbit_r27_c217 bl_217 br_217 wl_27 vdd gnd cell_6t
Xbit_r28_c217 bl_217 br_217 wl_28 vdd gnd cell_6t
Xbit_r29_c217 bl_217 br_217 wl_29 vdd gnd cell_6t
Xbit_r30_c217 bl_217 br_217 wl_30 vdd gnd cell_6t
Xbit_r31_c217 bl_217 br_217 wl_31 vdd gnd cell_6t
Xbit_r32_c217 bl_217 br_217 wl_32 vdd gnd cell_6t
Xbit_r33_c217 bl_217 br_217 wl_33 vdd gnd cell_6t
Xbit_r34_c217 bl_217 br_217 wl_34 vdd gnd cell_6t
Xbit_r35_c217 bl_217 br_217 wl_35 vdd gnd cell_6t
Xbit_r36_c217 bl_217 br_217 wl_36 vdd gnd cell_6t
Xbit_r37_c217 bl_217 br_217 wl_37 vdd gnd cell_6t
Xbit_r38_c217 bl_217 br_217 wl_38 vdd gnd cell_6t
Xbit_r39_c217 bl_217 br_217 wl_39 vdd gnd cell_6t
Xbit_r40_c217 bl_217 br_217 wl_40 vdd gnd cell_6t
Xbit_r41_c217 bl_217 br_217 wl_41 vdd gnd cell_6t
Xbit_r42_c217 bl_217 br_217 wl_42 vdd gnd cell_6t
Xbit_r43_c217 bl_217 br_217 wl_43 vdd gnd cell_6t
Xbit_r44_c217 bl_217 br_217 wl_44 vdd gnd cell_6t
Xbit_r45_c217 bl_217 br_217 wl_45 vdd gnd cell_6t
Xbit_r46_c217 bl_217 br_217 wl_46 vdd gnd cell_6t
Xbit_r47_c217 bl_217 br_217 wl_47 vdd gnd cell_6t
Xbit_r48_c217 bl_217 br_217 wl_48 vdd gnd cell_6t
Xbit_r49_c217 bl_217 br_217 wl_49 vdd gnd cell_6t
Xbit_r50_c217 bl_217 br_217 wl_50 vdd gnd cell_6t
Xbit_r51_c217 bl_217 br_217 wl_51 vdd gnd cell_6t
Xbit_r52_c217 bl_217 br_217 wl_52 vdd gnd cell_6t
Xbit_r53_c217 bl_217 br_217 wl_53 vdd gnd cell_6t
Xbit_r54_c217 bl_217 br_217 wl_54 vdd gnd cell_6t
Xbit_r55_c217 bl_217 br_217 wl_55 vdd gnd cell_6t
Xbit_r56_c217 bl_217 br_217 wl_56 vdd gnd cell_6t
Xbit_r57_c217 bl_217 br_217 wl_57 vdd gnd cell_6t
Xbit_r58_c217 bl_217 br_217 wl_58 vdd gnd cell_6t
Xbit_r59_c217 bl_217 br_217 wl_59 vdd gnd cell_6t
Xbit_r60_c217 bl_217 br_217 wl_60 vdd gnd cell_6t
Xbit_r61_c217 bl_217 br_217 wl_61 vdd gnd cell_6t
Xbit_r62_c217 bl_217 br_217 wl_62 vdd gnd cell_6t
Xbit_r63_c217 bl_217 br_217 wl_63 vdd gnd cell_6t
Xbit_r64_c217 bl_217 br_217 wl_64 vdd gnd cell_6t
Xbit_r65_c217 bl_217 br_217 wl_65 vdd gnd cell_6t
Xbit_r66_c217 bl_217 br_217 wl_66 vdd gnd cell_6t
Xbit_r67_c217 bl_217 br_217 wl_67 vdd gnd cell_6t
Xbit_r68_c217 bl_217 br_217 wl_68 vdd gnd cell_6t
Xbit_r69_c217 bl_217 br_217 wl_69 vdd gnd cell_6t
Xbit_r70_c217 bl_217 br_217 wl_70 vdd gnd cell_6t
Xbit_r71_c217 bl_217 br_217 wl_71 vdd gnd cell_6t
Xbit_r72_c217 bl_217 br_217 wl_72 vdd gnd cell_6t
Xbit_r73_c217 bl_217 br_217 wl_73 vdd gnd cell_6t
Xbit_r74_c217 bl_217 br_217 wl_74 vdd gnd cell_6t
Xbit_r75_c217 bl_217 br_217 wl_75 vdd gnd cell_6t
Xbit_r76_c217 bl_217 br_217 wl_76 vdd gnd cell_6t
Xbit_r77_c217 bl_217 br_217 wl_77 vdd gnd cell_6t
Xbit_r78_c217 bl_217 br_217 wl_78 vdd gnd cell_6t
Xbit_r79_c217 bl_217 br_217 wl_79 vdd gnd cell_6t
Xbit_r80_c217 bl_217 br_217 wl_80 vdd gnd cell_6t
Xbit_r81_c217 bl_217 br_217 wl_81 vdd gnd cell_6t
Xbit_r82_c217 bl_217 br_217 wl_82 vdd gnd cell_6t
Xbit_r83_c217 bl_217 br_217 wl_83 vdd gnd cell_6t
Xbit_r84_c217 bl_217 br_217 wl_84 vdd gnd cell_6t
Xbit_r85_c217 bl_217 br_217 wl_85 vdd gnd cell_6t
Xbit_r86_c217 bl_217 br_217 wl_86 vdd gnd cell_6t
Xbit_r87_c217 bl_217 br_217 wl_87 vdd gnd cell_6t
Xbit_r88_c217 bl_217 br_217 wl_88 vdd gnd cell_6t
Xbit_r89_c217 bl_217 br_217 wl_89 vdd gnd cell_6t
Xbit_r90_c217 bl_217 br_217 wl_90 vdd gnd cell_6t
Xbit_r91_c217 bl_217 br_217 wl_91 vdd gnd cell_6t
Xbit_r92_c217 bl_217 br_217 wl_92 vdd gnd cell_6t
Xbit_r93_c217 bl_217 br_217 wl_93 vdd gnd cell_6t
Xbit_r94_c217 bl_217 br_217 wl_94 vdd gnd cell_6t
Xbit_r95_c217 bl_217 br_217 wl_95 vdd gnd cell_6t
Xbit_r96_c217 bl_217 br_217 wl_96 vdd gnd cell_6t
Xbit_r97_c217 bl_217 br_217 wl_97 vdd gnd cell_6t
Xbit_r98_c217 bl_217 br_217 wl_98 vdd gnd cell_6t
Xbit_r99_c217 bl_217 br_217 wl_99 vdd gnd cell_6t
Xbit_r100_c217 bl_217 br_217 wl_100 vdd gnd cell_6t
Xbit_r101_c217 bl_217 br_217 wl_101 vdd gnd cell_6t
Xbit_r102_c217 bl_217 br_217 wl_102 vdd gnd cell_6t
Xbit_r103_c217 bl_217 br_217 wl_103 vdd gnd cell_6t
Xbit_r104_c217 bl_217 br_217 wl_104 vdd gnd cell_6t
Xbit_r105_c217 bl_217 br_217 wl_105 vdd gnd cell_6t
Xbit_r106_c217 bl_217 br_217 wl_106 vdd gnd cell_6t
Xbit_r107_c217 bl_217 br_217 wl_107 vdd gnd cell_6t
Xbit_r108_c217 bl_217 br_217 wl_108 vdd gnd cell_6t
Xbit_r109_c217 bl_217 br_217 wl_109 vdd gnd cell_6t
Xbit_r110_c217 bl_217 br_217 wl_110 vdd gnd cell_6t
Xbit_r111_c217 bl_217 br_217 wl_111 vdd gnd cell_6t
Xbit_r112_c217 bl_217 br_217 wl_112 vdd gnd cell_6t
Xbit_r113_c217 bl_217 br_217 wl_113 vdd gnd cell_6t
Xbit_r114_c217 bl_217 br_217 wl_114 vdd gnd cell_6t
Xbit_r115_c217 bl_217 br_217 wl_115 vdd gnd cell_6t
Xbit_r116_c217 bl_217 br_217 wl_116 vdd gnd cell_6t
Xbit_r117_c217 bl_217 br_217 wl_117 vdd gnd cell_6t
Xbit_r118_c217 bl_217 br_217 wl_118 vdd gnd cell_6t
Xbit_r119_c217 bl_217 br_217 wl_119 vdd gnd cell_6t
Xbit_r120_c217 bl_217 br_217 wl_120 vdd gnd cell_6t
Xbit_r121_c217 bl_217 br_217 wl_121 vdd gnd cell_6t
Xbit_r122_c217 bl_217 br_217 wl_122 vdd gnd cell_6t
Xbit_r123_c217 bl_217 br_217 wl_123 vdd gnd cell_6t
Xbit_r124_c217 bl_217 br_217 wl_124 vdd gnd cell_6t
Xbit_r125_c217 bl_217 br_217 wl_125 vdd gnd cell_6t
Xbit_r126_c217 bl_217 br_217 wl_126 vdd gnd cell_6t
Xbit_r127_c217 bl_217 br_217 wl_127 vdd gnd cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd cell_6t
Xbit_r1_c218 bl_218 br_218 wl_1 vdd gnd cell_6t
Xbit_r2_c218 bl_218 br_218 wl_2 vdd gnd cell_6t
Xbit_r3_c218 bl_218 br_218 wl_3 vdd gnd cell_6t
Xbit_r4_c218 bl_218 br_218 wl_4 vdd gnd cell_6t
Xbit_r5_c218 bl_218 br_218 wl_5 vdd gnd cell_6t
Xbit_r6_c218 bl_218 br_218 wl_6 vdd gnd cell_6t
Xbit_r7_c218 bl_218 br_218 wl_7 vdd gnd cell_6t
Xbit_r8_c218 bl_218 br_218 wl_8 vdd gnd cell_6t
Xbit_r9_c218 bl_218 br_218 wl_9 vdd gnd cell_6t
Xbit_r10_c218 bl_218 br_218 wl_10 vdd gnd cell_6t
Xbit_r11_c218 bl_218 br_218 wl_11 vdd gnd cell_6t
Xbit_r12_c218 bl_218 br_218 wl_12 vdd gnd cell_6t
Xbit_r13_c218 bl_218 br_218 wl_13 vdd gnd cell_6t
Xbit_r14_c218 bl_218 br_218 wl_14 vdd gnd cell_6t
Xbit_r15_c218 bl_218 br_218 wl_15 vdd gnd cell_6t
Xbit_r16_c218 bl_218 br_218 wl_16 vdd gnd cell_6t
Xbit_r17_c218 bl_218 br_218 wl_17 vdd gnd cell_6t
Xbit_r18_c218 bl_218 br_218 wl_18 vdd gnd cell_6t
Xbit_r19_c218 bl_218 br_218 wl_19 vdd gnd cell_6t
Xbit_r20_c218 bl_218 br_218 wl_20 vdd gnd cell_6t
Xbit_r21_c218 bl_218 br_218 wl_21 vdd gnd cell_6t
Xbit_r22_c218 bl_218 br_218 wl_22 vdd gnd cell_6t
Xbit_r23_c218 bl_218 br_218 wl_23 vdd gnd cell_6t
Xbit_r24_c218 bl_218 br_218 wl_24 vdd gnd cell_6t
Xbit_r25_c218 bl_218 br_218 wl_25 vdd gnd cell_6t
Xbit_r26_c218 bl_218 br_218 wl_26 vdd gnd cell_6t
Xbit_r27_c218 bl_218 br_218 wl_27 vdd gnd cell_6t
Xbit_r28_c218 bl_218 br_218 wl_28 vdd gnd cell_6t
Xbit_r29_c218 bl_218 br_218 wl_29 vdd gnd cell_6t
Xbit_r30_c218 bl_218 br_218 wl_30 vdd gnd cell_6t
Xbit_r31_c218 bl_218 br_218 wl_31 vdd gnd cell_6t
Xbit_r32_c218 bl_218 br_218 wl_32 vdd gnd cell_6t
Xbit_r33_c218 bl_218 br_218 wl_33 vdd gnd cell_6t
Xbit_r34_c218 bl_218 br_218 wl_34 vdd gnd cell_6t
Xbit_r35_c218 bl_218 br_218 wl_35 vdd gnd cell_6t
Xbit_r36_c218 bl_218 br_218 wl_36 vdd gnd cell_6t
Xbit_r37_c218 bl_218 br_218 wl_37 vdd gnd cell_6t
Xbit_r38_c218 bl_218 br_218 wl_38 vdd gnd cell_6t
Xbit_r39_c218 bl_218 br_218 wl_39 vdd gnd cell_6t
Xbit_r40_c218 bl_218 br_218 wl_40 vdd gnd cell_6t
Xbit_r41_c218 bl_218 br_218 wl_41 vdd gnd cell_6t
Xbit_r42_c218 bl_218 br_218 wl_42 vdd gnd cell_6t
Xbit_r43_c218 bl_218 br_218 wl_43 vdd gnd cell_6t
Xbit_r44_c218 bl_218 br_218 wl_44 vdd gnd cell_6t
Xbit_r45_c218 bl_218 br_218 wl_45 vdd gnd cell_6t
Xbit_r46_c218 bl_218 br_218 wl_46 vdd gnd cell_6t
Xbit_r47_c218 bl_218 br_218 wl_47 vdd gnd cell_6t
Xbit_r48_c218 bl_218 br_218 wl_48 vdd gnd cell_6t
Xbit_r49_c218 bl_218 br_218 wl_49 vdd gnd cell_6t
Xbit_r50_c218 bl_218 br_218 wl_50 vdd gnd cell_6t
Xbit_r51_c218 bl_218 br_218 wl_51 vdd gnd cell_6t
Xbit_r52_c218 bl_218 br_218 wl_52 vdd gnd cell_6t
Xbit_r53_c218 bl_218 br_218 wl_53 vdd gnd cell_6t
Xbit_r54_c218 bl_218 br_218 wl_54 vdd gnd cell_6t
Xbit_r55_c218 bl_218 br_218 wl_55 vdd gnd cell_6t
Xbit_r56_c218 bl_218 br_218 wl_56 vdd gnd cell_6t
Xbit_r57_c218 bl_218 br_218 wl_57 vdd gnd cell_6t
Xbit_r58_c218 bl_218 br_218 wl_58 vdd gnd cell_6t
Xbit_r59_c218 bl_218 br_218 wl_59 vdd gnd cell_6t
Xbit_r60_c218 bl_218 br_218 wl_60 vdd gnd cell_6t
Xbit_r61_c218 bl_218 br_218 wl_61 vdd gnd cell_6t
Xbit_r62_c218 bl_218 br_218 wl_62 vdd gnd cell_6t
Xbit_r63_c218 bl_218 br_218 wl_63 vdd gnd cell_6t
Xbit_r64_c218 bl_218 br_218 wl_64 vdd gnd cell_6t
Xbit_r65_c218 bl_218 br_218 wl_65 vdd gnd cell_6t
Xbit_r66_c218 bl_218 br_218 wl_66 vdd gnd cell_6t
Xbit_r67_c218 bl_218 br_218 wl_67 vdd gnd cell_6t
Xbit_r68_c218 bl_218 br_218 wl_68 vdd gnd cell_6t
Xbit_r69_c218 bl_218 br_218 wl_69 vdd gnd cell_6t
Xbit_r70_c218 bl_218 br_218 wl_70 vdd gnd cell_6t
Xbit_r71_c218 bl_218 br_218 wl_71 vdd gnd cell_6t
Xbit_r72_c218 bl_218 br_218 wl_72 vdd gnd cell_6t
Xbit_r73_c218 bl_218 br_218 wl_73 vdd gnd cell_6t
Xbit_r74_c218 bl_218 br_218 wl_74 vdd gnd cell_6t
Xbit_r75_c218 bl_218 br_218 wl_75 vdd gnd cell_6t
Xbit_r76_c218 bl_218 br_218 wl_76 vdd gnd cell_6t
Xbit_r77_c218 bl_218 br_218 wl_77 vdd gnd cell_6t
Xbit_r78_c218 bl_218 br_218 wl_78 vdd gnd cell_6t
Xbit_r79_c218 bl_218 br_218 wl_79 vdd gnd cell_6t
Xbit_r80_c218 bl_218 br_218 wl_80 vdd gnd cell_6t
Xbit_r81_c218 bl_218 br_218 wl_81 vdd gnd cell_6t
Xbit_r82_c218 bl_218 br_218 wl_82 vdd gnd cell_6t
Xbit_r83_c218 bl_218 br_218 wl_83 vdd gnd cell_6t
Xbit_r84_c218 bl_218 br_218 wl_84 vdd gnd cell_6t
Xbit_r85_c218 bl_218 br_218 wl_85 vdd gnd cell_6t
Xbit_r86_c218 bl_218 br_218 wl_86 vdd gnd cell_6t
Xbit_r87_c218 bl_218 br_218 wl_87 vdd gnd cell_6t
Xbit_r88_c218 bl_218 br_218 wl_88 vdd gnd cell_6t
Xbit_r89_c218 bl_218 br_218 wl_89 vdd gnd cell_6t
Xbit_r90_c218 bl_218 br_218 wl_90 vdd gnd cell_6t
Xbit_r91_c218 bl_218 br_218 wl_91 vdd gnd cell_6t
Xbit_r92_c218 bl_218 br_218 wl_92 vdd gnd cell_6t
Xbit_r93_c218 bl_218 br_218 wl_93 vdd gnd cell_6t
Xbit_r94_c218 bl_218 br_218 wl_94 vdd gnd cell_6t
Xbit_r95_c218 bl_218 br_218 wl_95 vdd gnd cell_6t
Xbit_r96_c218 bl_218 br_218 wl_96 vdd gnd cell_6t
Xbit_r97_c218 bl_218 br_218 wl_97 vdd gnd cell_6t
Xbit_r98_c218 bl_218 br_218 wl_98 vdd gnd cell_6t
Xbit_r99_c218 bl_218 br_218 wl_99 vdd gnd cell_6t
Xbit_r100_c218 bl_218 br_218 wl_100 vdd gnd cell_6t
Xbit_r101_c218 bl_218 br_218 wl_101 vdd gnd cell_6t
Xbit_r102_c218 bl_218 br_218 wl_102 vdd gnd cell_6t
Xbit_r103_c218 bl_218 br_218 wl_103 vdd gnd cell_6t
Xbit_r104_c218 bl_218 br_218 wl_104 vdd gnd cell_6t
Xbit_r105_c218 bl_218 br_218 wl_105 vdd gnd cell_6t
Xbit_r106_c218 bl_218 br_218 wl_106 vdd gnd cell_6t
Xbit_r107_c218 bl_218 br_218 wl_107 vdd gnd cell_6t
Xbit_r108_c218 bl_218 br_218 wl_108 vdd gnd cell_6t
Xbit_r109_c218 bl_218 br_218 wl_109 vdd gnd cell_6t
Xbit_r110_c218 bl_218 br_218 wl_110 vdd gnd cell_6t
Xbit_r111_c218 bl_218 br_218 wl_111 vdd gnd cell_6t
Xbit_r112_c218 bl_218 br_218 wl_112 vdd gnd cell_6t
Xbit_r113_c218 bl_218 br_218 wl_113 vdd gnd cell_6t
Xbit_r114_c218 bl_218 br_218 wl_114 vdd gnd cell_6t
Xbit_r115_c218 bl_218 br_218 wl_115 vdd gnd cell_6t
Xbit_r116_c218 bl_218 br_218 wl_116 vdd gnd cell_6t
Xbit_r117_c218 bl_218 br_218 wl_117 vdd gnd cell_6t
Xbit_r118_c218 bl_218 br_218 wl_118 vdd gnd cell_6t
Xbit_r119_c218 bl_218 br_218 wl_119 vdd gnd cell_6t
Xbit_r120_c218 bl_218 br_218 wl_120 vdd gnd cell_6t
Xbit_r121_c218 bl_218 br_218 wl_121 vdd gnd cell_6t
Xbit_r122_c218 bl_218 br_218 wl_122 vdd gnd cell_6t
Xbit_r123_c218 bl_218 br_218 wl_123 vdd gnd cell_6t
Xbit_r124_c218 bl_218 br_218 wl_124 vdd gnd cell_6t
Xbit_r125_c218 bl_218 br_218 wl_125 vdd gnd cell_6t
Xbit_r126_c218 bl_218 br_218 wl_126 vdd gnd cell_6t
Xbit_r127_c218 bl_218 br_218 wl_127 vdd gnd cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd cell_6t
Xbit_r1_c219 bl_219 br_219 wl_1 vdd gnd cell_6t
Xbit_r2_c219 bl_219 br_219 wl_2 vdd gnd cell_6t
Xbit_r3_c219 bl_219 br_219 wl_3 vdd gnd cell_6t
Xbit_r4_c219 bl_219 br_219 wl_4 vdd gnd cell_6t
Xbit_r5_c219 bl_219 br_219 wl_5 vdd gnd cell_6t
Xbit_r6_c219 bl_219 br_219 wl_6 vdd gnd cell_6t
Xbit_r7_c219 bl_219 br_219 wl_7 vdd gnd cell_6t
Xbit_r8_c219 bl_219 br_219 wl_8 vdd gnd cell_6t
Xbit_r9_c219 bl_219 br_219 wl_9 vdd gnd cell_6t
Xbit_r10_c219 bl_219 br_219 wl_10 vdd gnd cell_6t
Xbit_r11_c219 bl_219 br_219 wl_11 vdd gnd cell_6t
Xbit_r12_c219 bl_219 br_219 wl_12 vdd gnd cell_6t
Xbit_r13_c219 bl_219 br_219 wl_13 vdd gnd cell_6t
Xbit_r14_c219 bl_219 br_219 wl_14 vdd gnd cell_6t
Xbit_r15_c219 bl_219 br_219 wl_15 vdd gnd cell_6t
Xbit_r16_c219 bl_219 br_219 wl_16 vdd gnd cell_6t
Xbit_r17_c219 bl_219 br_219 wl_17 vdd gnd cell_6t
Xbit_r18_c219 bl_219 br_219 wl_18 vdd gnd cell_6t
Xbit_r19_c219 bl_219 br_219 wl_19 vdd gnd cell_6t
Xbit_r20_c219 bl_219 br_219 wl_20 vdd gnd cell_6t
Xbit_r21_c219 bl_219 br_219 wl_21 vdd gnd cell_6t
Xbit_r22_c219 bl_219 br_219 wl_22 vdd gnd cell_6t
Xbit_r23_c219 bl_219 br_219 wl_23 vdd gnd cell_6t
Xbit_r24_c219 bl_219 br_219 wl_24 vdd gnd cell_6t
Xbit_r25_c219 bl_219 br_219 wl_25 vdd gnd cell_6t
Xbit_r26_c219 bl_219 br_219 wl_26 vdd gnd cell_6t
Xbit_r27_c219 bl_219 br_219 wl_27 vdd gnd cell_6t
Xbit_r28_c219 bl_219 br_219 wl_28 vdd gnd cell_6t
Xbit_r29_c219 bl_219 br_219 wl_29 vdd gnd cell_6t
Xbit_r30_c219 bl_219 br_219 wl_30 vdd gnd cell_6t
Xbit_r31_c219 bl_219 br_219 wl_31 vdd gnd cell_6t
Xbit_r32_c219 bl_219 br_219 wl_32 vdd gnd cell_6t
Xbit_r33_c219 bl_219 br_219 wl_33 vdd gnd cell_6t
Xbit_r34_c219 bl_219 br_219 wl_34 vdd gnd cell_6t
Xbit_r35_c219 bl_219 br_219 wl_35 vdd gnd cell_6t
Xbit_r36_c219 bl_219 br_219 wl_36 vdd gnd cell_6t
Xbit_r37_c219 bl_219 br_219 wl_37 vdd gnd cell_6t
Xbit_r38_c219 bl_219 br_219 wl_38 vdd gnd cell_6t
Xbit_r39_c219 bl_219 br_219 wl_39 vdd gnd cell_6t
Xbit_r40_c219 bl_219 br_219 wl_40 vdd gnd cell_6t
Xbit_r41_c219 bl_219 br_219 wl_41 vdd gnd cell_6t
Xbit_r42_c219 bl_219 br_219 wl_42 vdd gnd cell_6t
Xbit_r43_c219 bl_219 br_219 wl_43 vdd gnd cell_6t
Xbit_r44_c219 bl_219 br_219 wl_44 vdd gnd cell_6t
Xbit_r45_c219 bl_219 br_219 wl_45 vdd gnd cell_6t
Xbit_r46_c219 bl_219 br_219 wl_46 vdd gnd cell_6t
Xbit_r47_c219 bl_219 br_219 wl_47 vdd gnd cell_6t
Xbit_r48_c219 bl_219 br_219 wl_48 vdd gnd cell_6t
Xbit_r49_c219 bl_219 br_219 wl_49 vdd gnd cell_6t
Xbit_r50_c219 bl_219 br_219 wl_50 vdd gnd cell_6t
Xbit_r51_c219 bl_219 br_219 wl_51 vdd gnd cell_6t
Xbit_r52_c219 bl_219 br_219 wl_52 vdd gnd cell_6t
Xbit_r53_c219 bl_219 br_219 wl_53 vdd gnd cell_6t
Xbit_r54_c219 bl_219 br_219 wl_54 vdd gnd cell_6t
Xbit_r55_c219 bl_219 br_219 wl_55 vdd gnd cell_6t
Xbit_r56_c219 bl_219 br_219 wl_56 vdd gnd cell_6t
Xbit_r57_c219 bl_219 br_219 wl_57 vdd gnd cell_6t
Xbit_r58_c219 bl_219 br_219 wl_58 vdd gnd cell_6t
Xbit_r59_c219 bl_219 br_219 wl_59 vdd gnd cell_6t
Xbit_r60_c219 bl_219 br_219 wl_60 vdd gnd cell_6t
Xbit_r61_c219 bl_219 br_219 wl_61 vdd gnd cell_6t
Xbit_r62_c219 bl_219 br_219 wl_62 vdd gnd cell_6t
Xbit_r63_c219 bl_219 br_219 wl_63 vdd gnd cell_6t
Xbit_r64_c219 bl_219 br_219 wl_64 vdd gnd cell_6t
Xbit_r65_c219 bl_219 br_219 wl_65 vdd gnd cell_6t
Xbit_r66_c219 bl_219 br_219 wl_66 vdd gnd cell_6t
Xbit_r67_c219 bl_219 br_219 wl_67 vdd gnd cell_6t
Xbit_r68_c219 bl_219 br_219 wl_68 vdd gnd cell_6t
Xbit_r69_c219 bl_219 br_219 wl_69 vdd gnd cell_6t
Xbit_r70_c219 bl_219 br_219 wl_70 vdd gnd cell_6t
Xbit_r71_c219 bl_219 br_219 wl_71 vdd gnd cell_6t
Xbit_r72_c219 bl_219 br_219 wl_72 vdd gnd cell_6t
Xbit_r73_c219 bl_219 br_219 wl_73 vdd gnd cell_6t
Xbit_r74_c219 bl_219 br_219 wl_74 vdd gnd cell_6t
Xbit_r75_c219 bl_219 br_219 wl_75 vdd gnd cell_6t
Xbit_r76_c219 bl_219 br_219 wl_76 vdd gnd cell_6t
Xbit_r77_c219 bl_219 br_219 wl_77 vdd gnd cell_6t
Xbit_r78_c219 bl_219 br_219 wl_78 vdd gnd cell_6t
Xbit_r79_c219 bl_219 br_219 wl_79 vdd gnd cell_6t
Xbit_r80_c219 bl_219 br_219 wl_80 vdd gnd cell_6t
Xbit_r81_c219 bl_219 br_219 wl_81 vdd gnd cell_6t
Xbit_r82_c219 bl_219 br_219 wl_82 vdd gnd cell_6t
Xbit_r83_c219 bl_219 br_219 wl_83 vdd gnd cell_6t
Xbit_r84_c219 bl_219 br_219 wl_84 vdd gnd cell_6t
Xbit_r85_c219 bl_219 br_219 wl_85 vdd gnd cell_6t
Xbit_r86_c219 bl_219 br_219 wl_86 vdd gnd cell_6t
Xbit_r87_c219 bl_219 br_219 wl_87 vdd gnd cell_6t
Xbit_r88_c219 bl_219 br_219 wl_88 vdd gnd cell_6t
Xbit_r89_c219 bl_219 br_219 wl_89 vdd gnd cell_6t
Xbit_r90_c219 bl_219 br_219 wl_90 vdd gnd cell_6t
Xbit_r91_c219 bl_219 br_219 wl_91 vdd gnd cell_6t
Xbit_r92_c219 bl_219 br_219 wl_92 vdd gnd cell_6t
Xbit_r93_c219 bl_219 br_219 wl_93 vdd gnd cell_6t
Xbit_r94_c219 bl_219 br_219 wl_94 vdd gnd cell_6t
Xbit_r95_c219 bl_219 br_219 wl_95 vdd gnd cell_6t
Xbit_r96_c219 bl_219 br_219 wl_96 vdd gnd cell_6t
Xbit_r97_c219 bl_219 br_219 wl_97 vdd gnd cell_6t
Xbit_r98_c219 bl_219 br_219 wl_98 vdd gnd cell_6t
Xbit_r99_c219 bl_219 br_219 wl_99 vdd gnd cell_6t
Xbit_r100_c219 bl_219 br_219 wl_100 vdd gnd cell_6t
Xbit_r101_c219 bl_219 br_219 wl_101 vdd gnd cell_6t
Xbit_r102_c219 bl_219 br_219 wl_102 vdd gnd cell_6t
Xbit_r103_c219 bl_219 br_219 wl_103 vdd gnd cell_6t
Xbit_r104_c219 bl_219 br_219 wl_104 vdd gnd cell_6t
Xbit_r105_c219 bl_219 br_219 wl_105 vdd gnd cell_6t
Xbit_r106_c219 bl_219 br_219 wl_106 vdd gnd cell_6t
Xbit_r107_c219 bl_219 br_219 wl_107 vdd gnd cell_6t
Xbit_r108_c219 bl_219 br_219 wl_108 vdd gnd cell_6t
Xbit_r109_c219 bl_219 br_219 wl_109 vdd gnd cell_6t
Xbit_r110_c219 bl_219 br_219 wl_110 vdd gnd cell_6t
Xbit_r111_c219 bl_219 br_219 wl_111 vdd gnd cell_6t
Xbit_r112_c219 bl_219 br_219 wl_112 vdd gnd cell_6t
Xbit_r113_c219 bl_219 br_219 wl_113 vdd gnd cell_6t
Xbit_r114_c219 bl_219 br_219 wl_114 vdd gnd cell_6t
Xbit_r115_c219 bl_219 br_219 wl_115 vdd gnd cell_6t
Xbit_r116_c219 bl_219 br_219 wl_116 vdd gnd cell_6t
Xbit_r117_c219 bl_219 br_219 wl_117 vdd gnd cell_6t
Xbit_r118_c219 bl_219 br_219 wl_118 vdd gnd cell_6t
Xbit_r119_c219 bl_219 br_219 wl_119 vdd gnd cell_6t
Xbit_r120_c219 bl_219 br_219 wl_120 vdd gnd cell_6t
Xbit_r121_c219 bl_219 br_219 wl_121 vdd gnd cell_6t
Xbit_r122_c219 bl_219 br_219 wl_122 vdd gnd cell_6t
Xbit_r123_c219 bl_219 br_219 wl_123 vdd gnd cell_6t
Xbit_r124_c219 bl_219 br_219 wl_124 vdd gnd cell_6t
Xbit_r125_c219 bl_219 br_219 wl_125 vdd gnd cell_6t
Xbit_r126_c219 bl_219 br_219 wl_126 vdd gnd cell_6t
Xbit_r127_c219 bl_219 br_219 wl_127 vdd gnd cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd cell_6t
Xbit_r1_c220 bl_220 br_220 wl_1 vdd gnd cell_6t
Xbit_r2_c220 bl_220 br_220 wl_2 vdd gnd cell_6t
Xbit_r3_c220 bl_220 br_220 wl_3 vdd gnd cell_6t
Xbit_r4_c220 bl_220 br_220 wl_4 vdd gnd cell_6t
Xbit_r5_c220 bl_220 br_220 wl_5 vdd gnd cell_6t
Xbit_r6_c220 bl_220 br_220 wl_6 vdd gnd cell_6t
Xbit_r7_c220 bl_220 br_220 wl_7 vdd gnd cell_6t
Xbit_r8_c220 bl_220 br_220 wl_8 vdd gnd cell_6t
Xbit_r9_c220 bl_220 br_220 wl_9 vdd gnd cell_6t
Xbit_r10_c220 bl_220 br_220 wl_10 vdd gnd cell_6t
Xbit_r11_c220 bl_220 br_220 wl_11 vdd gnd cell_6t
Xbit_r12_c220 bl_220 br_220 wl_12 vdd gnd cell_6t
Xbit_r13_c220 bl_220 br_220 wl_13 vdd gnd cell_6t
Xbit_r14_c220 bl_220 br_220 wl_14 vdd gnd cell_6t
Xbit_r15_c220 bl_220 br_220 wl_15 vdd gnd cell_6t
Xbit_r16_c220 bl_220 br_220 wl_16 vdd gnd cell_6t
Xbit_r17_c220 bl_220 br_220 wl_17 vdd gnd cell_6t
Xbit_r18_c220 bl_220 br_220 wl_18 vdd gnd cell_6t
Xbit_r19_c220 bl_220 br_220 wl_19 vdd gnd cell_6t
Xbit_r20_c220 bl_220 br_220 wl_20 vdd gnd cell_6t
Xbit_r21_c220 bl_220 br_220 wl_21 vdd gnd cell_6t
Xbit_r22_c220 bl_220 br_220 wl_22 vdd gnd cell_6t
Xbit_r23_c220 bl_220 br_220 wl_23 vdd gnd cell_6t
Xbit_r24_c220 bl_220 br_220 wl_24 vdd gnd cell_6t
Xbit_r25_c220 bl_220 br_220 wl_25 vdd gnd cell_6t
Xbit_r26_c220 bl_220 br_220 wl_26 vdd gnd cell_6t
Xbit_r27_c220 bl_220 br_220 wl_27 vdd gnd cell_6t
Xbit_r28_c220 bl_220 br_220 wl_28 vdd gnd cell_6t
Xbit_r29_c220 bl_220 br_220 wl_29 vdd gnd cell_6t
Xbit_r30_c220 bl_220 br_220 wl_30 vdd gnd cell_6t
Xbit_r31_c220 bl_220 br_220 wl_31 vdd gnd cell_6t
Xbit_r32_c220 bl_220 br_220 wl_32 vdd gnd cell_6t
Xbit_r33_c220 bl_220 br_220 wl_33 vdd gnd cell_6t
Xbit_r34_c220 bl_220 br_220 wl_34 vdd gnd cell_6t
Xbit_r35_c220 bl_220 br_220 wl_35 vdd gnd cell_6t
Xbit_r36_c220 bl_220 br_220 wl_36 vdd gnd cell_6t
Xbit_r37_c220 bl_220 br_220 wl_37 vdd gnd cell_6t
Xbit_r38_c220 bl_220 br_220 wl_38 vdd gnd cell_6t
Xbit_r39_c220 bl_220 br_220 wl_39 vdd gnd cell_6t
Xbit_r40_c220 bl_220 br_220 wl_40 vdd gnd cell_6t
Xbit_r41_c220 bl_220 br_220 wl_41 vdd gnd cell_6t
Xbit_r42_c220 bl_220 br_220 wl_42 vdd gnd cell_6t
Xbit_r43_c220 bl_220 br_220 wl_43 vdd gnd cell_6t
Xbit_r44_c220 bl_220 br_220 wl_44 vdd gnd cell_6t
Xbit_r45_c220 bl_220 br_220 wl_45 vdd gnd cell_6t
Xbit_r46_c220 bl_220 br_220 wl_46 vdd gnd cell_6t
Xbit_r47_c220 bl_220 br_220 wl_47 vdd gnd cell_6t
Xbit_r48_c220 bl_220 br_220 wl_48 vdd gnd cell_6t
Xbit_r49_c220 bl_220 br_220 wl_49 vdd gnd cell_6t
Xbit_r50_c220 bl_220 br_220 wl_50 vdd gnd cell_6t
Xbit_r51_c220 bl_220 br_220 wl_51 vdd gnd cell_6t
Xbit_r52_c220 bl_220 br_220 wl_52 vdd gnd cell_6t
Xbit_r53_c220 bl_220 br_220 wl_53 vdd gnd cell_6t
Xbit_r54_c220 bl_220 br_220 wl_54 vdd gnd cell_6t
Xbit_r55_c220 bl_220 br_220 wl_55 vdd gnd cell_6t
Xbit_r56_c220 bl_220 br_220 wl_56 vdd gnd cell_6t
Xbit_r57_c220 bl_220 br_220 wl_57 vdd gnd cell_6t
Xbit_r58_c220 bl_220 br_220 wl_58 vdd gnd cell_6t
Xbit_r59_c220 bl_220 br_220 wl_59 vdd gnd cell_6t
Xbit_r60_c220 bl_220 br_220 wl_60 vdd gnd cell_6t
Xbit_r61_c220 bl_220 br_220 wl_61 vdd gnd cell_6t
Xbit_r62_c220 bl_220 br_220 wl_62 vdd gnd cell_6t
Xbit_r63_c220 bl_220 br_220 wl_63 vdd gnd cell_6t
Xbit_r64_c220 bl_220 br_220 wl_64 vdd gnd cell_6t
Xbit_r65_c220 bl_220 br_220 wl_65 vdd gnd cell_6t
Xbit_r66_c220 bl_220 br_220 wl_66 vdd gnd cell_6t
Xbit_r67_c220 bl_220 br_220 wl_67 vdd gnd cell_6t
Xbit_r68_c220 bl_220 br_220 wl_68 vdd gnd cell_6t
Xbit_r69_c220 bl_220 br_220 wl_69 vdd gnd cell_6t
Xbit_r70_c220 bl_220 br_220 wl_70 vdd gnd cell_6t
Xbit_r71_c220 bl_220 br_220 wl_71 vdd gnd cell_6t
Xbit_r72_c220 bl_220 br_220 wl_72 vdd gnd cell_6t
Xbit_r73_c220 bl_220 br_220 wl_73 vdd gnd cell_6t
Xbit_r74_c220 bl_220 br_220 wl_74 vdd gnd cell_6t
Xbit_r75_c220 bl_220 br_220 wl_75 vdd gnd cell_6t
Xbit_r76_c220 bl_220 br_220 wl_76 vdd gnd cell_6t
Xbit_r77_c220 bl_220 br_220 wl_77 vdd gnd cell_6t
Xbit_r78_c220 bl_220 br_220 wl_78 vdd gnd cell_6t
Xbit_r79_c220 bl_220 br_220 wl_79 vdd gnd cell_6t
Xbit_r80_c220 bl_220 br_220 wl_80 vdd gnd cell_6t
Xbit_r81_c220 bl_220 br_220 wl_81 vdd gnd cell_6t
Xbit_r82_c220 bl_220 br_220 wl_82 vdd gnd cell_6t
Xbit_r83_c220 bl_220 br_220 wl_83 vdd gnd cell_6t
Xbit_r84_c220 bl_220 br_220 wl_84 vdd gnd cell_6t
Xbit_r85_c220 bl_220 br_220 wl_85 vdd gnd cell_6t
Xbit_r86_c220 bl_220 br_220 wl_86 vdd gnd cell_6t
Xbit_r87_c220 bl_220 br_220 wl_87 vdd gnd cell_6t
Xbit_r88_c220 bl_220 br_220 wl_88 vdd gnd cell_6t
Xbit_r89_c220 bl_220 br_220 wl_89 vdd gnd cell_6t
Xbit_r90_c220 bl_220 br_220 wl_90 vdd gnd cell_6t
Xbit_r91_c220 bl_220 br_220 wl_91 vdd gnd cell_6t
Xbit_r92_c220 bl_220 br_220 wl_92 vdd gnd cell_6t
Xbit_r93_c220 bl_220 br_220 wl_93 vdd gnd cell_6t
Xbit_r94_c220 bl_220 br_220 wl_94 vdd gnd cell_6t
Xbit_r95_c220 bl_220 br_220 wl_95 vdd gnd cell_6t
Xbit_r96_c220 bl_220 br_220 wl_96 vdd gnd cell_6t
Xbit_r97_c220 bl_220 br_220 wl_97 vdd gnd cell_6t
Xbit_r98_c220 bl_220 br_220 wl_98 vdd gnd cell_6t
Xbit_r99_c220 bl_220 br_220 wl_99 vdd gnd cell_6t
Xbit_r100_c220 bl_220 br_220 wl_100 vdd gnd cell_6t
Xbit_r101_c220 bl_220 br_220 wl_101 vdd gnd cell_6t
Xbit_r102_c220 bl_220 br_220 wl_102 vdd gnd cell_6t
Xbit_r103_c220 bl_220 br_220 wl_103 vdd gnd cell_6t
Xbit_r104_c220 bl_220 br_220 wl_104 vdd gnd cell_6t
Xbit_r105_c220 bl_220 br_220 wl_105 vdd gnd cell_6t
Xbit_r106_c220 bl_220 br_220 wl_106 vdd gnd cell_6t
Xbit_r107_c220 bl_220 br_220 wl_107 vdd gnd cell_6t
Xbit_r108_c220 bl_220 br_220 wl_108 vdd gnd cell_6t
Xbit_r109_c220 bl_220 br_220 wl_109 vdd gnd cell_6t
Xbit_r110_c220 bl_220 br_220 wl_110 vdd gnd cell_6t
Xbit_r111_c220 bl_220 br_220 wl_111 vdd gnd cell_6t
Xbit_r112_c220 bl_220 br_220 wl_112 vdd gnd cell_6t
Xbit_r113_c220 bl_220 br_220 wl_113 vdd gnd cell_6t
Xbit_r114_c220 bl_220 br_220 wl_114 vdd gnd cell_6t
Xbit_r115_c220 bl_220 br_220 wl_115 vdd gnd cell_6t
Xbit_r116_c220 bl_220 br_220 wl_116 vdd gnd cell_6t
Xbit_r117_c220 bl_220 br_220 wl_117 vdd gnd cell_6t
Xbit_r118_c220 bl_220 br_220 wl_118 vdd gnd cell_6t
Xbit_r119_c220 bl_220 br_220 wl_119 vdd gnd cell_6t
Xbit_r120_c220 bl_220 br_220 wl_120 vdd gnd cell_6t
Xbit_r121_c220 bl_220 br_220 wl_121 vdd gnd cell_6t
Xbit_r122_c220 bl_220 br_220 wl_122 vdd gnd cell_6t
Xbit_r123_c220 bl_220 br_220 wl_123 vdd gnd cell_6t
Xbit_r124_c220 bl_220 br_220 wl_124 vdd gnd cell_6t
Xbit_r125_c220 bl_220 br_220 wl_125 vdd gnd cell_6t
Xbit_r126_c220 bl_220 br_220 wl_126 vdd gnd cell_6t
Xbit_r127_c220 bl_220 br_220 wl_127 vdd gnd cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd cell_6t
Xbit_r1_c221 bl_221 br_221 wl_1 vdd gnd cell_6t
Xbit_r2_c221 bl_221 br_221 wl_2 vdd gnd cell_6t
Xbit_r3_c221 bl_221 br_221 wl_3 vdd gnd cell_6t
Xbit_r4_c221 bl_221 br_221 wl_4 vdd gnd cell_6t
Xbit_r5_c221 bl_221 br_221 wl_5 vdd gnd cell_6t
Xbit_r6_c221 bl_221 br_221 wl_6 vdd gnd cell_6t
Xbit_r7_c221 bl_221 br_221 wl_7 vdd gnd cell_6t
Xbit_r8_c221 bl_221 br_221 wl_8 vdd gnd cell_6t
Xbit_r9_c221 bl_221 br_221 wl_9 vdd gnd cell_6t
Xbit_r10_c221 bl_221 br_221 wl_10 vdd gnd cell_6t
Xbit_r11_c221 bl_221 br_221 wl_11 vdd gnd cell_6t
Xbit_r12_c221 bl_221 br_221 wl_12 vdd gnd cell_6t
Xbit_r13_c221 bl_221 br_221 wl_13 vdd gnd cell_6t
Xbit_r14_c221 bl_221 br_221 wl_14 vdd gnd cell_6t
Xbit_r15_c221 bl_221 br_221 wl_15 vdd gnd cell_6t
Xbit_r16_c221 bl_221 br_221 wl_16 vdd gnd cell_6t
Xbit_r17_c221 bl_221 br_221 wl_17 vdd gnd cell_6t
Xbit_r18_c221 bl_221 br_221 wl_18 vdd gnd cell_6t
Xbit_r19_c221 bl_221 br_221 wl_19 vdd gnd cell_6t
Xbit_r20_c221 bl_221 br_221 wl_20 vdd gnd cell_6t
Xbit_r21_c221 bl_221 br_221 wl_21 vdd gnd cell_6t
Xbit_r22_c221 bl_221 br_221 wl_22 vdd gnd cell_6t
Xbit_r23_c221 bl_221 br_221 wl_23 vdd gnd cell_6t
Xbit_r24_c221 bl_221 br_221 wl_24 vdd gnd cell_6t
Xbit_r25_c221 bl_221 br_221 wl_25 vdd gnd cell_6t
Xbit_r26_c221 bl_221 br_221 wl_26 vdd gnd cell_6t
Xbit_r27_c221 bl_221 br_221 wl_27 vdd gnd cell_6t
Xbit_r28_c221 bl_221 br_221 wl_28 vdd gnd cell_6t
Xbit_r29_c221 bl_221 br_221 wl_29 vdd gnd cell_6t
Xbit_r30_c221 bl_221 br_221 wl_30 vdd gnd cell_6t
Xbit_r31_c221 bl_221 br_221 wl_31 vdd gnd cell_6t
Xbit_r32_c221 bl_221 br_221 wl_32 vdd gnd cell_6t
Xbit_r33_c221 bl_221 br_221 wl_33 vdd gnd cell_6t
Xbit_r34_c221 bl_221 br_221 wl_34 vdd gnd cell_6t
Xbit_r35_c221 bl_221 br_221 wl_35 vdd gnd cell_6t
Xbit_r36_c221 bl_221 br_221 wl_36 vdd gnd cell_6t
Xbit_r37_c221 bl_221 br_221 wl_37 vdd gnd cell_6t
Xbit_r38_c221 bl_221 br_221 wl_38 vdd gnd cell_6t
Xbit_r39_c221 bl_221 br_221 wl_39 vdd gnd cell_6t
Xbit_r40_c221 bl_221 br_221 wl_40 vdd gnd cell_6t
Xbit_r41_c221 bl_221 br_221 wl_41 vdd gnd cell_6t
Xbit_r42_c221 bl_221 br_221 wl_42 vdd gnd cell_6t
Xbit_r43_c221 bl_221 br_221 wl_43 vdd gnd cell_6t
Xbit_r44_c221 bl_221 br_221 wl_44 vdd gnd cell_6t
Xbit_r45_c221 bl_221 br_221 wl_45 vdd gnd cell_6t
Xbit_r46_c221 bl_221 br_221 wl_46 vdd gnd cell_6t
Xbit_r47_c221 bl_221 br_221 wl_47 vdd gnd cell_6t
Xbit_r48_c221 bl_221 br_221 wl_48 vdd gnd cell_6t
Xbit_r49_c221 bl_221 br_221 wl_49 vdd gnd cell_6t
Xbit_r50_c221 bl_221 br_221 wl_50 vdd gnd cell_6t
Xbit_r51_c221 bl_221 br_221 wl_51 vdd gnd cell_6t
Xbit_r52_c221 bl_221 br_221 wl_52 vdd gnd cell_6t
Xbit_r53_c221 bl_221 br_221 wl_53 vdd gnd cell_6t
Xbit_r54_c221 bl_221 br_221 wl_54 vdd gnd cell_6t
Xbit_r55_c221 bl_221 br_221 wl_55 vdd gnd cell_6t
Xbit_r56_c221 bl_221 br_221 wl_56 vdd gnd cell_6t
Xbit_r57_c221 bl_221 br_221 wl_57 vdd gnd cell_6t
Xbit_r58_c221 bl_221 br_221 wl_58 vdd gnd cell_6t
Xbit_r59_c221 bl_221 br_221 wl_59 vdd gnd cell_6t
Xbit_r60_c221 bl_221 br_221 wl_60 vdd gnd cell_6t
Xbit_r61_c221 bl_221 br_221 wl_61 vdd gnd cell_6t
Xbit_r62_c221 bl_221 br_221 wl_62 vdd gnd cell_6t
Xbit_r63_c221 bl_221 br_221 wl_63 vdd gnd cell_6t
Xbit_r64_c221 bl_221 br_221 wl_64 vdd gnd cell_6t
Xbit_r65_c221 bl_221 br_221 wl_65 vdd gnd cell_6t
Xbit_r66_c221 bl_221 br_221 wl_66 vdd gnd cell_6t
Xbit_r67_c221 bl_221 br_221 wl_67 vdd gnd cell_6t
Xbit_r68_c221 bl_221 br_221 wl_68 vdd gnd cell_6t
Xbit_r69_c221 bl_221 br_221 wl_69 vdd gnd cell_6t
Xbit_r70_c221 bl_221 br_221 wl_70 vdd gnd cell_6t
Xbit_r71_c221 bl_221 br_221 wl_71 vdd gnd cell_6t
Xbit_r72_c221 bl_221 br_221 wl_72 vdd gnd cell_6t
Xbit_r73_c221 bl_221 br_221 wl_73 vdd gnd cell_6t
Xbit_r74_c221 bl_221 br_221 wl_74 vdd gnd cell_6t
Xbit_r75_c221 bl_221 br_221 wl_75 vdd gnd cell_6t
Xbit_r76_c221 bl_221 br_221 wl_76 vdd gnd cell_6t
Xbit_r77_c221 bl_221 br_221 wl_77 vdd gnd cell_6t
Xbit_r78_c221 bl_221 br_221 wl_78 vdd gnd cell_6t
Xbit_r79_c221 bl_221 br_221 wl_79 vdd gnd cell_6t
Xbit_r80_c221 bl_221 br_221 wl_80 vdd gnd cell_6t
Xbit_r81_c221 bl_221 br_221 wl_81 vdd gnd cell_6t
Xbit_r82_c221 bl_221 br_221 wl_82 vdd gnd cell_6t
Xbit_r83_c221 bl_221 br_221 wl_83 vdd gnd cell_6t
Xbit_r84_c221 bl_221 br_221 wl_84 vdd gnd cell_6t
Xbit_r85_c221 bl_221 br_221 wl_85 vdd gnd cell_6t
Xbit_r86_c221 bl_221 br_221 wl_86 vdd gnd cell_6t
Xbit_r87_c221 bl_221 br_221 wl_87 vdd gnd cell_6t
Xbit_r88_c221 bl_221 br_221 wl_88 vdd gnd cell_6t
Xbit_r89_c221 bl_221 br_221 wl_89 vdd gnd cell_6t
Xbit_r90_c221 bl_221 br_221 wl_90 vdd gnd cell_6t
Xbit_r91_c221 bl_221 br_221 wl_91 vdd gnd cell_6t
Xbit_r92_c221 bl_221 br_221 wl_92 vdd gnd cell_6t
Xbit_r93_c221 bl_221 br_221 wl_93 vdd gnd cell_6t
Xbit_r94_c221 bl_221 br_221 wl_94 vdd gnd cell_6t
Xbit_r95_c221 bl_221 br_221 wl_95 vdd gnd cell_6t
Xbit_r96_c221 bl_221 br_221 wl_96 vdd gnd cell_6t
Xbit_r97_c221 bl_221 br_221 wl_97 vdd gnd cell_6t
Xbit_r98_c221 bl_221 br_221 wl_98 vdd gnd cell_6t
Xbit_r99_c221 bl_221 br_221 wl_99 vdd gnd cell_6t
Xbit_r100_c221 bl_221 br_221 wl_100 vdd gnd cell_6t
Xbit_r101_c221 bl_221 br_221 wl_101 vdd gnd cell_6t
Xbit_r102_c221 bl_221 br_221 wl_102 vdd gnd cell_6t
Xbit_r103_c221 bl_221 br_221 wl_103 vdd gnd cell_6t
Xbit_r104_c221 bl_221 br_221 wl_104 vdd gnd cell_6t
Xbit_r105_c221 bl_221 br_221 wl_105 vdd gnd cell_6t
Xbit_r106_c221 bl_221 br_221 wl_106 vdd gnd cell_6t
Xbit_r107_c221 bl_221 br_221 wl_107 vdd gnd cell_6t
Xbit_r108_c221 bl_221 br_221 wl_108 vdd gnd cell_6t
Xbit_r109_c221 bl_221 br_221 wl_109 vdd gnd cell_6t
Xbit_r110_c221 bl_221 br_221 wl_110 vdd gnd cell_6t
Xbit_r111_c221 bl_221 br_221 wl_111 vdd gnd cell_6t
Xbit_r112_c221 bl_221 br_221 wl_112 vdd gnd cell_6t
Xbit_r113_c221 bl_221 br_221 wl_113 vdd gnd cell_6t
Xbit_r114_c221 bl_221 br_221 wl_114 vdd gnd cell_6t
Xbit_r115_c221 bl_221 br_221 wl_115 vdd gnd cell_6t
Xbit_r116_c221 bl_221 br_221 wl_116 vdd gnd cell_6t
Xbit_r117_c221 bl_221 br_221 wl_117 vdd gnd cell_6t
Xbit_r118_c221 bl_221 br_221 wl_118 vdd gnd cell_6t
Xbit_r119_c221 bl_221 br_221 wl_119 vdd gnd cell_6t
Xbit_r120_c221 bl_221 br_221 wl_120 vdd gnd cell_6t
Xbit_r121_c221 bl_221 br_221 wl_121 vdd gnd cell_6t
Xbit_r122_c221 bl_221 br_221 wl_122 vdd gnd cell_6t
Xbit_r123_c221 bl_221 br_221 wl_123 vdd gnd cell_6t
Xbit_r124_c221 bl_221 br_221 wl_124 vdd gnd cell_6t
Xbit_r125_c221 bl_221 br_221 wl_125 vdd gnd cell_6t
Xbit_r126_c221 bl_221 br_221 wl_126 vdd gnd cell_6t
Xbit_r127_c221 bl_221 br_221 wl_127 vdd gnd cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd cell_6t
Xbit_r1_c222 bl_222 br_222 wl_1 vdd gnd cell_6t
Xbit_r2_c222 bl_222 br_222 wl_2 vdd gnd cell_6t
Xbit_r3_c222 bl_222 br_222 wl_3 vdd gnd cell_6t
Xbit_r4_c222 bl_222 br_222 wl_4 vdd gnd cell_6t
Xbit_r5_c222 bl_222 br_222 wl_5 vdd gnd cell_6t
Xbit_r6_c222 bl_222 br_222 wl_6 vdd gnd cell_6t
Xbit_r7_c222 bl_222 br_222 wl_7 vdd gnd cell_6t
Xbit_r8_c222 bl_222 br_222 wl_8 vdd gnd cell_6t
Xbit_r9_c222 bl_222 br_222 wl_9 vdd gnd cell_6t
Xbit_r10_c222 bl_222 br_222 wl_10 vdd gnd cell_6t
Xbit_r11_c222 bl_222 br_222 wl_11 vdd gnd cell_6t
Xbit_r12_c222 bl_222 br_222 wl_12 vdd gnd cell_6t
Xbit_r13_c222 bl_222 br_222 wl_13 vdd gnd cell_6t
Xbit_r14_c222 bl_222 br_222 wl_14 vdd gnd cell_6t
Xbit_r15_c222 bl_222 br_222 wl_15 vdd gnd cell_6t
Xbit_r16_c222 bl_222 br_222 wl_16 vdd gnd cell_6t
Xbit_r17_c222 bl_222 br_222 wl_17 vdd gnd cell_6t
Xbit_r18_c222 bl_222 br_222 wl_18 vdd gnd cell_6t
Xbit_r19_c222 bl_222 br_222 wl_19 vdd gnd cell_6t
Xbit_r20_c222 bl_222 br_222 wl_20 vdd gnd cell_6t
Xbit_r21_c222 bl_222 br_222 wl_21 vdd gnd cell_6t
Xbit_r22_c222 bl_222 br_222 wl_22 vdd gnd cell_6t
Xbit_r23_c222 bl_222 br_222 wl_23 vdd gnd cell_6t
Xbit_r24_c222 bl_222 br_222 wl_24 vdd gnd cell_6t
Xbit_r25_c222 bl_222 br_222 wl_25 vdd gnd cell_6t
Xbit_r26_c222 bl_222 br_222 wl_26 vdd gnd cell_6t
Xbit_r27_c222 bl_222 br_222 wl_27 vdd gnd cell_6t
Xbit_r28_c222 bl_222 br_222 wl_28 vdd gnd cell_6t
Xbit_r29_c222 bl_222 br_222 wl_29 vdd gnd cell_6t
Xbit_r30_c222 bl_222 br_222 wl_30 vdd gnd cell_6t
Xbit_r31_c222 bl_222 br_222 wl_31 vdd gnd cell_6t
Xbit_r32_c222 bl_222 br_222 wl_32 vdd gnd cell_6t
Xbit_r33_c222 bl_222 br_222 wl_33 vdd gnd cell_6t
Xbit_r34_c222 bl_222 br_222 wl_34 vdd gnd cell_6t
Xbit_r35_c222 bl_222 br_222 wl_35 vdd gnd cell_6t
Xbit_r36_c222 bl_222 br_222 wl_36 vdd gnd cell_6t
Xbit_r37_c222 bl_222 br_222 wl_37 vdd gnd cell_6t
Xbit_r38_c222 bl_222 br_222 wl_38 vdd gnd cell_6t
Xbit_r39_c222 bl_222 br_222 wl_39 vdd gnd cell_6t
Xbit_r40_c222 bl_222 br_222 wl_40 vdd gnd cell_6t
Xbit_r41_c222 bl_222 br_222 wl_41 vdd gnd cell_6t
Xbit_r42_c222 bl_222 br_222 wl_42 vdd gnd cell_6t
Xbit_r43_c222 bl_222 br_222 wl_43 vdd gnd cell_6t
Xbit_r44_c222 bl_222 br_222 wl_44 vdd gnd cell_6t
Xbit_r45_c222 bl_222 br_222 wl_45 vdd gnd cell_6t
Xbit_r46_c222 bl_222 br_222 wl_46 vdd gnd cell_6t
Xbit_r47_c222 bl_222 br_222 wl_47 vdd gnd cell_6t
Xbit_r48_c222 bl_222 br_222 wl_48 vdd gnd cell_6t
Xbit_r49_c222 bl_222 br_222 wl_49 vdd gnd cell_6t
Xbit_r50_c222 bl_222 br_222 wl_50 vdd gnd cell_6t
Xbit_r51_c222 bl_222 br_222 wl_51 vdd gnd cell_6t
Xbit_r52_c222 bl_222 br_222 wl_52 vdd gnd cell_6t
Xbit_r53_c222 bl_222 br_222 wl_53 vdd gnd cell_6t
Xbit_r54_c222 bl_222 br_222 wl_54 vdd gnd cell_6t
Xbit_r55_c222 bl_222 br_222 wl_55 vdd gnd cell_6t
Xbit_r56_c222 bl_222 br_222 wl_56 vdd gnd cell_6t
Xbit_r57_c222 bl_222 br_222 wl_57 vdd gnd cell_6t
Xbit_r58_c222 bl_222 br_222 wl_58 vdd gnd cell_6t
Xbit_r59_c222 bl_222 br_222 wl_59 vdd gnd cell_6t
Xbit_r60_c222 bl_222 br_222 wl_60 vdd gnd cell_6t
Xbit_r61_c222 bl_222 br_222 wl_61 vdd gnd cell_6t
Xbit_r62_c222 bl_222 br_222 wl_62 vdd gnd cell_6t
Xbit_r63_c222 bl_222 br_222 wl_63 vdd gnd cell_6t
Xbit_r64_c222 bl_222 br_222 wl_64 vdd gnd cell_6t
Xbit_r65_c222 bl_222 br_222 wl_65 vdd gnd cell_6t
Xbit_r66_c222 bl_222 br_222 wl_66 vdd gnd cell_6t
Xbit_r67_c222 bl_222 br_222 wl_67 vdd gnd cell_6t
Xbit_r68_c222 bl_222 br_222 wl_68 vdd gnd cell_6t
Xbit_r69_c222 bl_222 br_222 wl_69 vdd gnd cell_6t
Xbit_r70_c222 bl_222 br_222 wl_70 vdd gnd cell_6t
Xbit_r71_c222 bl_222 br_222 wl_71 vdd gnd cell_6t
Xbit_r72_c222 bl_222 br_222 wl_72 vdd gnd cell_6t
Xbit_r73_c222 bl_222 br_222 wl_73 vdd gnd cell_6t
Xbit_r74_c222 bl_222 br_222 wl_74 vdd gnd cell_6t
Xbit_r75_c222 bl_222 br_222 wl_75 vdd gnd cell_6t
Xbit_r76_c222 bl_222 br_222 wl_76 vdd gnd cell_6t
Xbit_r77_c222 bl_222 br_222 wl_77 vdd gnd cell_6t
Xbit_r78_c222 bl_222 br_222 wl_78 vdd gnd cell_6t
Xbit_r79_c222 bl_222 br_222 wl_79 vdd gnd cell_6t
Xbit_r80_c222 bl_222 br_222 wl_80 vdd gnd cell_6t
Xbit_r81_c222 bl_222 br_222 wl_81 vdd gnd cell_6t
Xbit_r82_c222 bl_222 br_222 wl_82 vdd gnd cell_6t
Xbit_r83_c222 bl_222 br_222 wl_83 vdd gnd cell_6t
Xbit_r84_c222 bl_222 br_222 wl_84 vdd gnd cell_6t
Xbit_r85_c222 bl_222 br_222 wl_85 vdd gnd cell_6t
Xbit_r86_c222 bl_222 br_222 wl_86 vdd gnd cell_6t
Xbit_r87_c222 bl_222 br_222 wl_87 vdd gnd cell_6t
Xbit_r88_c222 bl_222 br_222 wl_88 vdd gnd cell_6t
Xbit_r89_c222 bl_222 br_222 wl_89 vdd gnd cell_6t
Xbit_r90_c222 bl_222 br_222 wl_90 vdd gnd cell_6t
Xbit_r91_c222 bl_222 br_222 wl_91 vdd gnd cell_6t
Xbit_r92_c222 bl_222 br_222 wl_92 vdd gnd cell_6t
Xbit_r93_c222 bl_222 br_222 wl_93 vdd gnd cell_6t
Xbit_r94_c222 bl_222 br_222 wl_94 vdd gnd cell_6t
Xbit_r95_c222 bl_222 br_222 wl_95 vdd gnd cell_6t
Xbit_r96_c222 bl_222 br_222 wl_96 vdd gnd cell_6t
Xbit_r97_c222 bl_222 br_222 wl_97 vdd gnd cell_6t
Xbit_r98_c222 bl_222 br_222 wl_98 vdd gnd cell_6t
Xbit_r99_c222 bl_222 br_222 wl_99 vdd gnd cell_6t
Xbit_r100_c222 bl_222 br_222 wl_100 vdd gnd cell_6t
Xbit_r101_c222 bl_222 br_222 wl_101 vdd gnd cell_6t
Xbit_r102_c222 bl_222 br_222 wl_102 vdd gnd cell_6t
Xbit_r103_c222 bl_222 br_222 wl_103 vdd gnd cell_6t
Xbit_r104_c222 bl_222 br_222 wl_104 vdd gnd cell_6t
Xbit_r105_c222 bl_222 br_222 wl_105 vdd gnd cell_6t
Xbit_r106_c222 bl_222 br_222 wl_106 vdd gnd cell_6t
Xbit_r107_c222 bl_222 br_222 wl_107 vdd gnd cell_6t
Xbit_r108_c222 bl_222 br_222 wl_108 vdd gnd cell_6t
Xbit_r109_c222 bl_222 br_222 wl_109 vdd gnd cell_6t
Xbit_r110_c222 bl_222 br_222 wl_110 vdd gnd cell_6t
Xbit_r111_c222 bl_222 br_222 wl_111 vdd gnd cell_6t
Xbit_r112_c222 bl_222 br_222 wl_112 vdd gnd cell_6t
Xbit_r113_c222 bl_222 br_222 wl_113 vdd gnd cell_6t
Xbit_r114_c222 bl_222 br_222 wl_114 vdd gnd cell_6t
Xbit_r115_c222 bl_222 br_222 wl_115 vdd gnd cell_6t
Xbit_r116_c222 bl_222 br_222 wl_116 vdd gnd cell_6t
Xbit_r117_c222 bl_222 br_222 wl_117 vdd gnd cell_6t
Xbit_r118_c222 bl_222 br_222 wl_118 vdd gnd cell_6t
Xbit_r119_c222 bl_222 br_222 wl_119 vdd gnd cell_6t
Xbit_r120_c222 bl_222 br_222 wl_120 vdd gnd cell_6t
Xbit_r121_c222 bl_222 br_222 wl_121 vdd gnd cell_6t
Xbit_r122_c222 bl_222 br_222 wl_122 vdd gnd cell_6t
Xbit_r123_c222 bl_222 br_222 wl_123 vdd gnd cell_6t
Xbit_r124_c222 bl_222 br_222 wl_124 vdd gnd cell_6t
Xbit_r125_c222 bl_222 br_222 wl_125 vdd gnd cell_6t
Xbit_r126_c222 bl_222 br_222 wl_126 vdd gnd cell_6t
Xbit_r127_c222 bl_222 br_222 wl_127 vdd gnd cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd cell_6t
Xbit_r1_c223 bl_223 br_223 wl_1 vdd gnd cell_6t
Xbit_r2_c223 bl_223 br_223 wl_2 vdd gnd cell_6t
Xbit_r3_c223 bl_223 br_223 wl_3 vdd gnd cell_6t
Xbit_r4_c223 bl_223 br_223 wl_4 vdd gnd cell_6t
Xbit_r5_c223 bl_223 br_223 wl_5 vdd gnd cell_6t
Xbit_r6_c223 bl_223 br_223 wl_6 vdd gnd cell_6t
Xbit_r7_c223 bl_223 br_223 wl_7 vdd gnd cell_6t
Xbit_r8_c223 bl_223 br_223 wl_8 vdd gnd cell_6t
Xbit_r9_c223 bl_223 br_223 wl_9 vdd gnd cell_6t
Xbit_r10_c223 bl_223 br_223 wl_10 vdd gnd cell_6t
Xbit_r11_c223 bl_223 br_223 wl_11 vdd gnd cell_6t
Xbit_r12_c223 bl_223 br_223 wl_12 vdd gnd cell_6t
Xbit_r13_c223 bl_223 br_223 wl_13 vdd gnd cell_6t
Xbit_r14_c223 bl_223 br_223 wl_14 vdd gnd cell_6t
Xbit_r15_c223 bl_223 br_223 wl_15 vdd gnd cell_6t
Xbit_r16_c223 bl_223 br_223 wl_16 vdd gnd cell_6t
Xbit_r17_c223 bl_223 br_223 wl_17 vdd gnd cell_6t
Xbit_r18_c223 bl_223 br_223 wl_18 vdd gnd cell_6t
Xbit_r19_c223 bl_223 br_223 wl_19 vdd gnd cell_6t
Xbit_r20_c223 bl_223 br_223 wl_20 vdd gnd cell_6t
Xbit_r21_c223 bl_223 br_223 wl_21 vdd gnd cell_6t
Xbit_r22_c223 bl_223 br_223 wl_22 vdd gnd cell_6t
Xbit_r23_c223 bl_223 br_223 wl_23 vdd gnd cell_6t
Xbit_r24_c223 bl_223 br_223 wl_24 vdd gnd cell_6t
Xbit_r25_c223 bl_223 br_223 wl_25 vdd gnd cell_6t
Xbit_r26_c223 bl_223 br_223 wl_26 vdd gnd cell_6t
Xbit_r27_c223 bl_223 br_223 wl_27 vdd gnd cell_6t
Xbit_r28_c223 bl_223 br_223 wl_28 vdd gnd cell_6t
Xbit_r29_c223 bl_223 br_223 wl_29 vdd gnd cell_6t
Xbit_r30_c223 bl_223 br_223 wl_30 vdd gnd cell_6t
Xbit_r31_c223 bl_223 br_223 wl_31 vdd gnd cell_6t
Xbit_r32_c223 bl_223 br_223 wl_32 vdd gnd cell_6t
Xbit_r33_c223 bl_223 br_223 wl_33 vdd gnd cell_6t
Xbit_r34_c223 bl_223 br_223 wl_34 vdd gnd cell_6t
Xbit_r35_c223 bl_223 br_223 wl_35 vdd gnd cell_6t
Xbit_r36_c223 bl_223 br_223 wl_36 vdd gnd cell_6t
Xbit_r37_c223 bl_223 br_223 wl_37 vdd gnd cell_6t
Xbit_r38_c223 bl_223 br_223 wl_38 vdd gnd cell_6t
Xbit_r39_c223 bl_223 br_223 wl_39 vdd gnd cell_6t
Xbit_r40_c223 bl_223 br_223 wl_40 vdd gnd cell_6t
Xbit_r41_c223 bl_223 br_223 wl_41 vdd gnd cell_6t
Xbit_r42_c223 bl_223 br_223 wl_42 vdd gnd cell_6t
Xbit_r43_c223 bl_223 br_223 wl_43 vdd gnd cell_6t
Xbit_r44_c223 bl_223 br_223 wl_44 vdd gnd cell_6t
Xbit_r45_c223 bl_223 br_223 wl_45 vdd gnd cell_6t
Xbit_r46_c223 bl_223 br_223 wl_46 vdd gnd cell_6t
Xbit_r47_c223 bl_223 br_223 wl_47 vdd gnd cell_6t
Xbit_r48_c223 bl_223 br_223 wl_48 vdd gnd cell_6t
Xbit_r49_c223 bl_223 br_223 wl_49 vdd gnd cell_6t
Xbit_r50_c223 bl_223 br_223 wl_50 vdd gnd cell_6t
Xbit_r51_c223 bl_223 br_223 wl_51 vdd gnd cell_6t
Xbit_r52_c223 bl_223 br_223 wl_52 vdd gnd cell_6t
Xbit_r53_c223 bl_223 br_223 wl_53 vdd gnd cell_6t
Xbit_r54_c223 bl_223 br_223 wl_54 vdd gnd cell_6t
Xbit_r55_c223 bl_223 br_223 wl_55 vdd gnd cell_6t
Xbit_r56_c223 bl_223 br_223 wl_56 vdd gnd cell_6t
Xbit_r57_c223 bl_223 br_223 wl_57 vdd gnd cell_6t
Xbit_r58_c223 bl_223 br_223 wl_58 vdd gnd cell_6t
Xbit_r59_c223 bl_223 br_223 wl_59 vdd gnd cell_6t
Xbit_r60_c223 bl_223 br_223 wl_60 vdd gnd cell_6t
Xbit_r61_c223 bl_223 br_223 wl_61 vdd gnd cell_6t
Xbit_r62_c223 bl_223 br_223 wl_62 vdd gnd cell_6t
Xbit_r63_c223 bl_223 br_223 wl_63 vdd gnd cell_6t
Xbit_r64_c223 bl_223 br_223 wl_64 vdd gnd cell_6t
Xbit_r65_c223 bl_223 br_223 wl_65 vdd gnd cell_6t
Xbit_r66_c223 bl_223 br_223 wl_66 vdd gnd cell_6t
Xbit_r67_c223 bl_223 br_223 wl_67 vdd gnd cell_6t
Xbit_r68_c223 bl_223 br_223 wl_68 vdd gnd cell_6t
Xbit_r69_c223 bl_223 br_223 wl_69 vdd gnd cell_6t
Xbit_r70_c223 bl_223 br_223 wl_70 vdd gnd cell_6t
Xbit_r71_c223 bl_223 br_223 wl_71 vdd gnd cell_6t
Xbit_r72_c223 bl_223 br_223 wl_72 vdd gnd cell_6t
Xbit_r73_c223 bl_223 br_223 wl_73 vdd gnd cell_6t
Xbit_r74_c223 bl_223 br_223 wl_74 vdd gnd cell_6t
Xbit_r75_c223 bl_223 br_223 wl_75 vdd gnd cell_6t
Xbit_r76_c223 bl_223 br_223 wl_76 vdd gnd cell_6t
Xbit_r77_c223 bl_223 br_223 wl_77 vdd gnd cell_6t
Xbit_r78_c223 bl_223 br_223 wl_78 vdd gnd cell_6t
Xbit_r79_c223 bl_223 br_223 wl_79 vdd gnd cell_6t
Xbit_r80_c223 bl_223 br_223 wl_80 vdd gnd cell_6t
Xbit_r81_c223 bl_223 br_223 wl_81 vdd gnd cell_6t
Xbit_r82_c223 bl_223 br_223 wl_82 vdd gnd cell_6t
Xbit_r83_c223 bl_223 br_223 wl_83 vdd gnd cell_6t
Xbit_r84_c223 bl_223 br_223 wl_84 vdd gnd cell_6t
Xbit_r85_c223 bl_223 br_223 wl_85 vdd gnd cell_6t
Xbit_r86_c223 bl_223 br_223 wl_86 vdd gnd cell_6t
Xbit_r87_c223 bl_223 br_223 wl_87 vdd gnd cell_6t
Xbit_r88_c223 bl_223 br_223 wl_88 vdd gnd cell_6t
Xbit_r89_c223 bl_223 br_223 wl_89 vdd gnd cell_6t
Xbit_r90_c223 bl_223 br_223 wl_90 vdd gnd cell_6t
Xbit_r91_c223 bl_223 br_223 wl_91 vdd gnd cell_6t
Xbit_r92_c223 bl_223 br_223 wl_92 vdd gnd cell_6t
Xbit_r93_c223 bl_223 br_223 wl_93 vdd gnd cell_6t
Xbit_r94_c223 bl_223 br_223 wl_94 vdd gnd cell_6t
Xbit_r95_c223 bl_223 br_223 wl_95 vdd gnd cell_6t
Xbit_r96_c223 bl_223 br_223 wl_96 vdd gnd cell_6t
Xbit_r97_c223 bl_223 br_223 wl_97 vdd gnd cell_6t
Xbit_r98_c223 bl_223 br_223 wl_98 vdd gnd cell_6t
Xbit_r99_c223 bl_223 br_223 wl_99 vdd gnd cell_6t
Xbit_r100_c223 bl_223 br_223 wl_100 vdd gnd cell_6t
Xbit_r101_c223 bl_223 br_223 wl_101 vdd gnd cell_6t
Xbit_r102_c223 bl_223 br_223 wl_102 vdd gnd cell_6t
Xbit_r103_c223 bl_223 br_223 wl_103 vdd gnd cell_6t
Xbit_r104_c223 bl_223 br_223 wl_104 vdd gnd cell_6t
Xbit_r105_c223 bl_223 br_223 wl_105 vdd gnd cell_6t
Xbit_r106_c223 bl_223 br_223 wl_106 vdd gnd cell_6t
Xbit_r107_c223 bl_223 br_223 wl_107 vdd gnd cell_6t
Xbit_r108_c223 bl_223 br_223 wl_108 vdd gnd cell_6t
Xbit_r109_c223 bl_223 br_223 wl_109 vdd gnd cell_6t
Xbit_r110_c223 bl_223 br_223 wl_110 vdd gnd cell_6t
Xbit_r111_c223 bl_223 br_223 wl_111 vdd gnd cell_6t
Xbit_r112_c223 bl_223 br_223 wl_112 vdd gnd cell_6t
Xbit_r113_c223 bl_223 br_223 wl_113 vdd gnd cell_6t
Xbit_r114_c223 bl_223 br_223 wl_114 vdd gnd cell_6t
Xbit_r115_c223 bl_223 br_223 wl_115 vdd gnd cell_6t
Xbit_r116_c223 bl_223 br_223 wl_116 vdd gnd cell_6t
Xbit_r117_c223 bl_223 br_223 wl_117 vdd gnd cell_6t
Xbit_r118_c223 bl_223 br_223 wl_118 vdd gnd cell_6t
Xbit_r119_c223 bl_223 br_223 wl_119 vdd gnd cell_6t
Xbit_r120_c223 bl_223 br_223 wl_120 vdd gnd cell_6t
Xbit_r121_c223 bl_223 br_223 wl_121 vdd gnd cell_6t
Xbit_r122_c223 bl_223 br_223 wl_122 vdd gnd cell_6t
Xbit_r123_c223 bl_223 br_223 wl_123 vdd gnd cell_6t
Xbit_r124_c223 bl_223 br_223 wl_124 vdd gnd cell_6t
Xbit_r125_c223 bl_223 br_223 wl_125 vdd gnd cell_6t
Xbit_r126_c223 bl_223 br_223 wl_126 vdd gnd cell_6t
Xbit_r127_c223 bl_223 br_223 wl_127 vdd gnd cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd cell_6t
Xbit_r1_c224 bl_224 br_224 wl_1 vdd gnd cell_6t
Xbit_r2_c224 bl_224 br_224 wl_2 vdd gnd cell_6t
Xbit_r3_c224 bl_224 br_224 wl_3 vdd gnd cell_6t
Xbit_r4_c224 bl_224 br_224 wl_4 vdd gnd cell_6t
Xbit_r5_c224 bl_224 br_224 wl_5 vdd gnd cell_6t
Xbit_r6_c224 bl_224 br_224 wl_6 vdd gnd cell_6t
Xbit_r7_c224 bl_224 br_224 wl_7 vdd gnd cell_6t
Xbit_r8_c224 bl_224 br_224 wl_8 vdd gnd cell_6t
Xbit_r9_c224 bl_224 br_224 wl_9 vdd gnd cell_6t
Xbit_r10_c224 bl_224 br_224 wl_10 vdd gnd cell_6t
Xbit_r11_c224 bl_224 br_224 wl_11 vdd gnd cell_6t
Xbit_r12_c224 bl_224 br_224 wl_12 vdd gnd cell_6t
Xbit_r13_c224 bl_224 br_224 wl_13 vdd gnd cell_6t
Xbit_r14_c224 bl_224 br_224 wl_14 vdd gnd cell_6t
Xbit_r15_c224 bl_224 br_224 wl_15 vdd gnd cell_6t
Xbit_r16_c224 bl_224 br_224 wl_16 vdd gnd cell_6t
Xbit_r17_c224 bl_224 br_224 wl_17 vdd gnd cell_6t
Xbit_r18_c224 bl_224 br_224 wl_18 vdd gnd cell_6t
Xbit_r19_c224 bl_224 br_224 wl_19 vdd gnd cell_6t
Xbit_r20_c224 bl_224 br_224 wl_20 vdd gnd cell_6t
Xbit_r21_c224 bl_224 br_224 wl_21 vdd gnd cell_6t
Xbit_r22_c224 bl_224 br_224 wl_22 vdd gnd cell_6t
Xbit_r23_c224 bl_224 br_224 wl_23 vdd gnd cell_6t
Xbit_r24_c224 bl_224 br_224 wl_24 vdd gnd cell_6t
Xbit_r25_c224 bl_224 br_224 wl_25 vdd gnd cell_6t
Xbit_r26_c224 bl_224 br_224 wl_26 vdd gnd cell_6t
Xbit_r27_c224 bl_224 br_224 wl_27 vdd gnd cell_6t
Xbit_r28_c224 bl_224 br_224 wl_28 vdd gnd cell_6t
Xbit_r29_c224 bl_224 br_224 wl_29 vdd gnd cell_6t
Xbit_r30_c224 bl_224 br_224 wl_30 vdd gnd cell_6t
Xbit_r31_c224 bl_224 br_224 wl_31 vdd gnd cell_6t
Xbit_r32_c224 bl_224 br_224 wl_32 vdd gnd cell_6t
Xbit_r33_c224 bl_224 br_224 wl_33 vdd gnd cell_6t
Xbit_r34_c224 bl_224 br_224 wl_34 vdd gnd cell_6t
Xbit_r35_c224 bl_224 br_224 wl_35 vdd gnd cell_6t
Xbit_r36_c224 bl_224 br_224 wl_36 vdd gnd cell_6t
Xbit_r37_c224 bl_224 br_224 wl_37 vdd gnd cell_6t
Xbit_r38_c224 bl_224 br_224 wl_38 vdd gnd cell_6t
Xbit_r39_c224 bl_224 br_224 wl_39 vdd gnd cell_6t
Xbit_r40_c224 bl_224 br_224 wl_40 vdd gnd cell_6t
Xbit_r41_c224 bl_224 br_224 wl_41 vdd gnd cell_6t
Xbit_r42_c224 bl_224 br_224 wl_42 vdd gnd cell_6t
Xbit_r43_c224 bl_224 br_224 wl_43 vdd gnd cell_6t
Xbit_r44_c224 bl_224 br_224 wl_44 vdd gnd cell_6t
Xbit_r45_c224 bl_224 br_224 wl_45 vdd gnd cell_6t
Xbit_r46_c224 bl_224 br_224 wl_46 vdd gnd cell_6t
Xbit_r47_c224 bl_224 br_224 wl_47 vdd gnd cell_6t
Xbit_r48_c224 bl_224 br_224 wl_48 vdd gnd cell_6t
Xbit_r49_c224 bl_224 br_224 wl_49 vdd gnd cell_6t
Xbit_r50_c224 bl_224 br_224 wl_50 vdd gnd cell_6t
Xbit_r51_c224 bl_224 br_224 wl_51 vdd gnd cell_6t
Xbit_r52_c224 bl_224 br_224 wl_52 vdd gnd cell_6t
Xbit_r53_c224 bl_224 br_224 wl_53 vdd gnd cell_6t
Xbit_r54_c224 bl_224 br_224 wl_54 vdd gnd cell_6t
Xbit_r55_c224 bl_224 br_224 wl_55 vdd gnd cell_6t
Xbit_r56_c224 bl_224 br_224 wl_56 vdd gnd cell_6t
Xbit_r57_c224 bl_224 br_224 wl_57 vdd gnd cell_6t
Xbit_r58_c224 bl_224 br_224 wl_58 vdd gnd cell_6t
Xbit_r59_c224 bl_224 br_224 wl_59 vdd gnd cell_6t
Xbit_r60_c224 bl_224 br_224 wl_60 vdd gnd cell_6t
Xbit_r61_c224 bl_224 br_224 wl_61 vdd gnd cell_6t
Xbit_r62_c224 bl_224 br_224 wl_62 vdd gnd cell_6t
Xbit_r63_c224 bl_224 br_224 wl_63 vdd gnd cell_6t
Xbit_r64_c224 bl_224 br_224 wl_64 vdd gnd cell_6t
Xbit_r65_c224 bl_224 br_224 wl_65 vdd gnd cell_6t
Xbit_r66_c224 bl_224 br_224 wl_66 vdd gnd cell_6t
Xbit_r67_c224 bl_224 br_224 wl_67 vdd gnd cell_6t
Xbit_r68_c224 bl_224 br_224 wl_68 vdd gnd cell_6t
Xbit_r69_c224 bl_224 br_224 wl_69 vdd gnd cell_6t
Xbit_r70_c224 bl_224 br_224 wl_70 vdd gnd cell_6t
Xbit_r71_c224 bl_224 br_224 wl_71 vdd gnd cell_6t
Xbit_r72_c224 bl_224 br_224 wl_72 vdd gnd cell_6t
Xbit_r73_c224 bl_224 br_224 wl_73 vdd gnd cell_6t
Xbit_r74_c224 bl_224 br_224 wl_74 vdd gnd cell_6t
Xbit_r75_c224 bl_224 br_224 wl_75 vdd gnd cell_6t
Xbit_r76_c224 bl_224 br_224 wl_76 vdd gnd cell_6t
Xbit_r77_c224 bl_224 br_224 wl_77 vdd gnd cell_6t
Xbit_r78_c224 bl_224 br_224 wl_78 vdd gnd cell_6t
Xbit_r79_c224 bl_224 br_224 wl_79 vdd gnd cell_6t
Xbit_r80_c224 bl_224 br_224 wl_80 vdd gnd cell_6t
Xbit_r81_c224 bl_224 br_224 wl_81 vdd gnd cell_6t
Xbit_r82_c224 bl_224 br_224 wl_82 vdd gnd cell_6t
Xbit_r83_c224 bl_224 br_224 wl_83 vdd gnd cell_6t
Xbit_r84_c224 bl_224 br_224 wl_84 vdd gnd cell_6t
Xbit_r85_c224 bl_224 br_224 wl_85 vdd gnd cell_6t
Xbit_r86_c224 bl_224 br_224 wl_86 vdd gnd cell_6t
Xbit_r87_c224 bl_224 br_224 wl_87 vdd gnd cell_6t
Xbit_r88_c224 bl_224 br_224 wl_88 vdd gnd cell_6t
Xbit_r89_c224 bl_224 br_224 wl_89 vdd gnd cell_6t
Xbit_r90_c224 bl_224 br_224 wl_90 vdd gnd cell_6t
Xbit_r91_c224 bl_224 br_224 wl_91 vdd gnd cell_6t
Xbit_r92_c224 bl_224 br_224 wl_92 vdd gnd cell_6t
Xbit_r93_c224 bl_224 br_224 wl_93 vdd gnd cell_6t
Xbit_r94_c224 bl_224 br_224 wl_94 vdd gnd cell_6t
Xbit_r95_c224 bl_224 br_224 wl_95 vdd gnd cell_6t
Xbit_r96_c224 bl_224 br_224 wl_96 vdd gnd cell_6t
Xbit_r97_c224 bl_224 br_224 wl_97 vdd gnd cell_6t
Xbit_r98_c224 bl_224 br_224 wl_98 vdd gnd cell_6t
Xbit_r99_c224 bl_224 br_224 wl_99 vdd gnd cell_6t
Xbit_r100_c224 bl_224 br_224 wl_100 vdd gnd cell_6t
Xbit_r101_c224 bl_224 br_224 wl_101 vdd gnd cell_6t
Xbit_r102_c224 bl_224 br_224 wl_102 vdd gnd cell_6t
Xbit_r103_c224 bl_224 br_224 wl_103 vdd gnd cell_6t
Xbit_r104_c224 bl_224 br_224 wl_104 vdd gnd cell_6t
Xbit_r105_c224 bl_224 br_224 wl_105 vdd gnd cell_6t
Xbit_r106_c224 bl_224 br_224 wl_106 vdd gnd cell_6t
Xbit_r107_c224 bl_224 br_224 wl_107 vdd gnd cell_6t
Xbit_r108_c224 bl_224 br_224 wl_108 vdd gnd cell_6t
Xbit_r109_c224 bl_224 br_224 wl_109 vdd gnd cell_6t
Xbit_r110_c224 bl_224 br_224 wl_110 vdd gnd cell_6t
Xbit_r111_c224 bl_224 br_224 wl_111 vdd gnd cell_6t
Xbit_r112_c224 bl_224 br_224 wl_112 vdd gnd cell_6t
Xbit_r113_c224 bl_224 br_224 wl_113 vdd gnd cell_6t
Xbit_r114_c224 bl_224 br_224 wl_114 vdd gnd cell_6t
Xbit_r115_c224 bl_224 br_224 wl_115 vdd gnd cell_6t
Xbit_r116_c224 bl_224 br_224 wl_116 vdd gnd cell_6t
Xbit_r117_c224 bl_224 br_224 wl_117 vdd gnd cell_6t
Xbit_r118_c224 bl_224 br_224 wl_118 vdd gnd cell_6t
Xbit_r119_c224 bl_224 br_224 wl_119 vdd gnd cell_6t
Xbit_r120_c224 bl_224 br_224 wl_120 vdd gnd cell_6t
Xbit_r121_c224 bl_224 br_224 wl_121 vdd gnd cell_6t
Xbit_r122_c224 bl_224 br_224 wl_122 vdd gnd cell_6t
Xbit_r123_c224 bl_224 br_224 wl_123 vdd gnd cell_6t
Xbit_r124_c224 bl_224 br_224 wl_124 vdd gnd cell_6t
Xbit_r125_c224 bl_224 br_224 wl_125 vdd gnd cell_6t
Xbit_r126_c224 bl_224 br_224 wl_126 vdd gnd cell_6t
Xbit_r127_c224 bl_224 br_224 wl_127 vdd gnd cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd cell_6t
Xbit_r1_c225 bl_225 br_225 wl_1 vdd gnd cell_6t
Xbit_r2_c225 bl_225 br_225 wl_2 vdd gnd cell_6t
Xbit_r3_c225 bl_225 br_225 wl_3 vdd gnd cell_6t
Xbit_r4_c225 bl_225 br_225 wl_4 vdd gnd cell_6t
Xbit_r5_c225 bl_225 br_225 wl_5 vdd gnd cell_6t
Xbit_r6_c225 bl_225 br_225 wl_6 vdd gnd cell_6t
Xbit_r7_c225 bl_225 br_225 wl_7 vdd gnd cell_6t
Xbit_r8_c225 bl_225 br_225 wl_8 vdd gnd cell_6t
Xbit_r9_c225 bl_225 br_225 wl_9 vdd gnd cell_6t
Xbit_r10_c225 bl_225 br_225 wl_10 vdd gnd cell_6t
Xbit_r11_c225 bl_225 br_225 wl_11 vdd gnd cell_6t
Xbit_r12_c225 bl_225 br_225 wl_12 vdd gnd cell_6t
Xbit_r13_c225 bl_225 br_225 wl_13 vdd gnd cell_6t
Xbit_r14_c225 bl_225 br_225 wl_14 vdd gnd cell_6t
Xbit_r15_c225 bl_225 br_225 wl_15 vdd gnd cell_6t
Xbit_r16_c225 bl_225 br_225 wl_16 vdd gnd cell_6t
Xbit_r17_c225 bl_225 br_225 wl_17 vdd gnd cell_6t
Xbit_r18_c225 bl_225 br_225 wl_18 vdd gnd cell_6t
Xbit_r19_c225 bl_225 br_225 wl_19 vdd gnd cell_6t
Xbit_r20_c225 bl_225 br_225 wl_20 vdd gnd cell_6t
Xbit_r21_c225 bl_225 br_225 wl_21 vdd gnd cell_6t
Xbit_r22_c225 bl_225 br_225 wl_22 vdd gnd cell_6t
Xbit_r23_c225 bl_225 br_225 wl_23 vdd gnd cell_6t
Xbit_r24_c225 bl_225 br_225 wl_24 vdd gnd cell_6t
Xbit_r25_c225 bl_225 br_225 wl_25 vdd gnd cell_6t
Xbit_r26_c225 bl_225 br_225 wl_26 vdd gnd cell_6t
Xbit_r27_c225 bl_225 br_225 wl_27 vdd gnd cell_6t
Xbit_r28_c225 bl_225 br_225 wl_28 vdd gnd cell_6t
Xbit_r29_c225 bl_225 br_225 wl_29 vdd gnd cell_6t
Xbit_r30_c225 bl_225 br_225 wl_30 vdd gnd cell_6t
Xbit_r31_c225 bl_225 br_225 wl_31 vdd gnd cell_6t
Xbit_r32_c225 bl_225 br_225 wl_32 vdd gnd cell_6t
Xbit_r33_c225 bl_225 br_225 wl_33 vdd gnd cell_6t
Xbit_r34_c225 bl_225 br_225 wl_34 vdd gnd cell_6t
Xbit_r35_c225 bl_225 br_225 wl_35 vdd gnd cell_6t
Xbit_r36_c225 bl_225 br_225 wl_36 vdd gnd cell_6t
Xbit_r37_c225 bl_225 br_225 wl_37 vdd gnd cell_6t
Xbit_r38_c225 bl_225 br_225 wl_38 vdd gnd cell_6t
Xbit_r39_c225 bl_225 br_225 wl_39 vdd gnd cell_6t
Xbit_r40_c225 bl_225 br_225 wl_40 vdd gnd cell_6t
Xbit_r41_c225 bl_225 br_225 wl_41 vdd gnd cell_6t
Xbit_r42_c225 bl_225 br_225 wl_42 vdd gnd cell_6t
Xbit_r43_c225 bl_225 br_225 wl_43 vdd gnd cell_6t
Xbit_r44_c225 bl_225 br_225 wl_44 vdd gnd cell_6t
Xbit_r45_c225 bl_225 br_225 wl_45 vdd gnd cell_6t
Xbit_r46_c225 bl_225 br_225 wl_46 vdd gnd cell_6t
Xbit_r47_c225 bl_225 br_225 wl_47 vdd gnd cell_6t
Xbit_r48_c225 bl_225 br_225 wl_48 vdd gnd cell_6t
Xbit_r49_c225 bl_225 br_225 wl_49 vdd gnd cell_6t
Xbit_r50_c225 bl_225 br_225 wl_50 vdd gnd cell_6t
Xbit_r51_c225 bl_225 br_225 wl_51 vdd gnd cell_6t
Xbit_r52_c225 bl_225 br_225 wl_52 vdd gnd cell_6t
Xbit_r53_c225 bl_225 br_225 wl_53 vdd gnd cell_6t
Xbit_r54_c225 bl_225 br_225 wl_54 vdd gnd cell_6t
Xbit_r55_c225 bl_225 br_225 wl_55 vdd gnd cell_6t
Xbit_r56_c225 bl_225 br_225 wl_56 vdd gnd cell_6t
Xbit_r57_c225 bl_225 br_225 wl_57 vdd gnd cell_6t
Xbit_r58_c225 bl_225 br_225 wl_58 vdd gnd cell_6t
Xbit_r59_c225 bl_225 br_225 wl_59 vdd gnd cell_6t
Xbit_r60_c225 bl_225 br_225 wl_60 vdd gnd cell_6t
Xbit_r61_c225 bl_225 br_225 wl_61 vdd gnd cell_6t
Xbit_r62_c225 bl_225 br_225 wl_62 vdd gnd cell_6t
Xbit_r63_c225 bl_225 br_225 wl_63 vdd gnd cell_6t
Xbit_r64_c225 bl_225 br_225 wl_64 vdd gnd cell_6t
Xbit_r65_c225 bl_225 br_225 wl_65 vdd gnd cell_6t
Xbit_r66_c225 bl_225 br_225 wl_66 vdd gnd cell_6t
Xbit_r67_c225 bl_225 br_225 wl_67 vdd gnd cell_6t
Xbit_r68_c225 bl_225 br_225 wl_68 vdd gnd cell_6t
Xbit_r69_c225 bl_225 br_225 wl_69 vdd gnd cell_6t
Xbit_r70_c225 bl_225 br_225 wl_70 vdd gnd cell_6t
Xbit_r71_c225 bl_225 br_225 wl_71 vdd gnd cell_6t
Xbit_r72_c225 bl_225 br_225 wl_72 vdd gnd cell_6t
Xbit_r73_c225 bl_225 br_225 wl_73 vdd gnd cell_6t
Xbit_r74_c225 bl_225 br_225 wl_74 vdd gnd cell_6t
Xbit_r75_c225 bl_225 br_225 wl_75 vdd gnd cell_6t
Xbit_r76_c225 bl_225 br_225 wl_76 vdd gnd cell_6t
Xbit_r77_c225 bl_225 br_225 wl_77 vdd gnd cell_6t
Xbit_r78_c225 bl_225 br_225 wl_78 vdd gnd cell_6t
Xbit_r79_c225 bl_225 br_225 wl_79 vdd gnd cell_6t
Xbit_r80_c225 bl_225 br_225 wl_80 vdd gnd cell_6t
Xbit_r81_c225 bl_225 br_225 wl_81 vdd gnd cell_6t
Xbit_r82_c225 bl_225 br_225 wl_82 vdd gnd cell_6t
Xbit_r83_c225 bl_225 br_225 wl_83 vdd gnd cell_6t
Xbit_r84_c225 bl_225 br_225 wl_84 vdd gnd cell_6t
Xbit_r85_c225 bl_225 br_225 wl_85 vdd gnd cell_6t
Xbit_r86_c225 bl_225 br_225 wl_86 vdd gnd cell_6t
Xbit_r87_c225 bl_225 br_225 wl_87 vdd gnd cell_6t
Xbit_r88_c225 bl_225 br_225 wl_88 vdd gnd cell_6t
Xbit_r89_c225 bl_225 br_225 wl_89 vdd gnd cell_6t
Xbit_r90_c225 bl_225 br_225 wl_90 vdd gnd cell_6t
Xbit_r91_c225 bl_225 br_225 wl_91 vdd gnd cell_6t
Xbit_r92_c225 bl_225 br_225 wl_92 vdd gnd cell_6t
Xbit_r93_c225 bl_225 br_225 wl_93 vdd gnd cell_6t
Xbit_r94_c225 bl_225 br_225 wl_94 vdd gnd cell_6t
Xbit_r95_c225 bl_225 br_225 wl_95 vdd gnd cell_6t
Xbit_r96_c225 bl_225 br_225 wl_96 vdd gnd cell_6t
Xbit_r97_c225 bl_225 br_225 wl_97 vdd gnd cell_6t
Xbit_r98_c225 bl_225 br_225 wl_98 vdd gnd cell_6t
Xbit_r99_c225 bl_225 br_225 wl_99 vdd gnd cell_6t
Xbit_r100_c225 bl_225 br_225 wl_100 vdd gnd cell_6t
Xbit_r101_c225 bl_225 br_225 wl_101 vdd gnd cell_6t
Xbit_r102_c225 bl_225 br_225 wl_102 vdd gnd cell_6t
Xbit_r103_c225 bl_225 br_225 wl_103 vdd gnd cell_6t
Xbit_r104_c225 bl_225 br_225 wl_104 vdd gnd cell_6t
Xbit_r105_c225 bl_225 br_225 wl_105 vdd gnd cell_6t
Xbit_r106_c225 bl_225 br_225 wl_106 vdd gnd cell_6t
Xbit_r107_c225 bl_225 br_225 wl_107 vdd gnd cell_6t
Xbit_r108_c225 bl_225 br_225 wl_108 vdd gnd cell_6t
Xbit_r109_c225 bl_225 br_225 wl_109 vdd gnd cell_6t
Xbit_r110_c225 bl_225 br_225 wl_110 vdd gnd cell_6t
Xbit_r111_c225 bl_225 br_225 wl_111 vdd gnd cell_6t
Xbit_r112_c225 bl_225 br_225 wl_112 vdd gnd cell_6t
Xbit_r113_c225 bl_225 br_225 wl_113 vdd gnd cell_6t
Xbit_r114_c225 bl_225 br_225 wl_114 vdd gnd cell_6t
Xbit_r115_c225 bl_225 br_225 wl_115 vdd gnd cell_6t
Xbit_r116_c225 bl_225 br_225 wl_116 vdd gnd cell_6t
Xbit_r117_c225 bl_225 br_225 wl_117 vdd gnd cell_6t
Xbit_r118_c225 bl_225 br_225 wl_118 vdd gnd cell_6t
Xbit_r119_c225 bl_225 br_225 wl_119 vdd gnd cell_6t
Xbit_r120_c225 bl_225 br_225 wl_120 vdd gnd cell_6t
Xbit_r121_c225 bl_225 br_225 wl_121 vdd gnd cell_6t
Xbit_r122_c225 bl_225 br_225 wl_122 vdd gnd cell_6t
Xbit_r123_c225 bl_225 br_225 wl_123 vdd gnd cell_6t
Xbit_r124_c225 bl_225 br_225 wl_124 vdd gnd cell_6t
Xbit_r125_c225 bl_225 br_225 wl_125 vdd gnd cell_6t
Xbit_r126_c225 bl_225 br_225 wl_126 vdd gnd cell_6t
Xbit_r127_c225 bl_225 br_225 wl_127 vdd gnd cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd cell_6t
Xbit_r1_c226 bl_226 br_226 wl_1 vdd gnd cell_6t
Xbit_r2_c226 bl_226 br_226 wl_2 vdd gnd cell_6t
Xbit_r3_c226 bl_226 br_226 wl_3 vdd gnd cell_6t
Xbit_r4_c226 bl_226 br_226 wl_4 vdd gnd cell_6t
Xbit_r5_c226 bl_226 br_226 wl_5 vdd gnd cell_6t
Xbit_r6_c226 bl_226 br_226 wl_6 vdd gnd cell_6t
Xbit_r7_c226 bl_226 br_226 wl_7 vdd gnd cell_6t
Xbit_r8_c226 bl_226 br_226 wl_8 vdd gnd cell_6t
Xbit_r9_c226 bl_226 br_226 wl_9 vdd gnd cell_6t
Xbit_r10_c226 bl_226 br_226 wl_10 vdd gnd cell_6t
Xbit_r11_c226 bl_226 br_226 wl_11 vdd gnd cell_6t
Xbit_r12_c226 bl_226 br_226 wl_12 vdd gnd cell_6t
Xbit_r13_c226 bl_226 br_226 wl_13 vdd gnd cell_6t
Xbit_r14_c226 bl_226 br_226 wl_14 vdd gnd cell_6t
Xbit_r15_c226 bl_226 br_226 wl_15 vdd gnd cell_6t
Xbit_r16_c226 bl_226 br_226 wl_16 vdd gnd cell_6t
Xbit_r17_c226 bl_226 br_226 wl_17 vdd gnd cell_6t
Xbit_r18_c226 bl_226 br_226 wl_18 vdd gnd cell_6t
Xbit_r19_c226 bl_226 br_226 wl_19 vdd gnd cell_6t
Xbit_r20_c226 bl_226 br_226 wl_20 vdd gnd cell_6t
Xbit_r21_c226 bl_226 br_226 wl_21 vdd gnd cell_6t
Xbit_r22_c226 bl_226 br_226 wl_22 vdd gnd cell_6t
Xbit_r23_c226 bl_226 br_226 wl_23 vdd gnd cell_6t
Xbit_r24_c226 bl_226 br_226 wl_24 vdd gnd cell_6t
Xbit_r25_c226 bl_226 br_226 wl_25 vdd gnd cell_6t
Xbit_r26_c226 bl_226 br_226 wl_26 vdd gnd cell_6t
Xbit_r27_c226 bl_226 br_226 wl_27 vdd gnd cell_6t
Xbit_r28_c226 bl_226 br_226 wl_28 vdd gnd cell_6t
Xbit_r29_c226 bl_226 br_226 wl_29 vdd gnd cell_6t
Xbit_r30_c226 bl_226 br_226 wl_30 vdd gnd cell_6t
Xbit_r31_c226 bl_226 br_226 wl_31 vdd gnd cell_6t
Xbit_r32_c226 bl_226 br_226 wl_32 vdd gnd cell_6t
Xbit_r33_c226 bl_226 br_226 wl_33 vdd gnd cell_6t
Xbit_r34_c226 bl_226 br_226 wl_34 vdd gnd cell_6t
Xbit_r35_c226 bl_226 br_226 wl_35 vdd gnd cell_6t
Xbit_r36_c226 bl_226 br_226 wl_36 vdd gnd cell_6t
Xbit_r37_c226 bl_226 br_226 wl_37 vdd gnd cell_6t
Xbit_r38_c226 bl_226 br_226 wl_38 vdd gnd cell_6t
Xbit_r39_c226 bl_226 br_226 wl_39 vdd gnd cell_6t
Xbit_r40_c226 bl_226 br_226 wl_40 vdd gnd cell_6t
Xbit_r41_c226 bl_226 br_226 wl_41 vdd gnd cell_6t
Xbit_r42_c226 bl_226 br_226 wl_42 vdd gnd cell_6t
Xbit_r43_c226 bl_226 br_226 wl_43 vdd gnd cell_6t
Xbit_r44_c226 bl_226 br_226 wl_44 vdd gnd cell_6t
Xbit_r45_c226 bl_226 br_226 wl_45 vdd gnd cell_6t
Xbit_r46_c226 bl_226 br_226 wl_46 vdd gnd cell_6t
Xbit_r47_c226 bl_226 br_226 wl_47 vdd gnd cell_6t
Xbit_r48_c226 bl_226 br_226 wl_48 vdd gnd cell_6t
Xbit_r49_c226 bl_226 br_226 wl_49 vdd gnd cell_6t
Xbit_r50_c226 bl_226 br_226 wl_50 vdd gnd cell_6t
Xbit_r51_c226 bl_226 br_226 wl_51 vdd gnd cell_6t
Xbit_r52_c226 bl_226 br_226 wl_52 vdd gnd cell_6t
Xbit_r53_c226 bl_226 br_226 wl_53 vdd gnd cell_6t
Xbit_r54_c226 bl_226 br_226 wl_54 vdd gnd cell_6t
Xbit_r55_c226 bl_226 br_226 wl_55 vdd gnd cell_6t
Xbit_r56_c226 bl_226 br_226 wl_56 vdd gnd cell_6t
Xbit_r57_c226 bl_226 br_226 wl_57 vdd gnd cell_6t
Xbit_r58_c226 bl_226 br_226 wl_58 vdd gnd cell_6t
Xbit_r59_c226 bl_226 br_226 wl_59 vdd gnd cell_6t
Xbit_r60_c226 bl_226 br_226 wl_60 vdd gnd cell_6t
Xbit_r61_c226 bl_226 br_226 wl_61 vdd gnd cell_6t
Xbit_r62_c226 bl_226 br_226 wl_62 vdd gnd cell_6t
Xbit_r63_c226 bl_226 br_226 wl_63 vdd gnd cell_6t
Xbit_r64_c226 bl_226 br_226 wl_64 vdd gnd cell_6t
Xbit_r65_c226 bl_226 br_226 wl_65 vdd gnd cell_6t
Xbit_r66_c226 bl_226 br_226 wl_66 vdd gnd cell_6t
Xbit_r67_c226 bl_226 br_226 wl_67 vdd gnd cell_6t
Xbit_r68_c226 bl_226 br_226 wl_68 vdd gnd cell_6t
Xbit_r69_c226 bl_226 br_226 wl_69 vdd gnd cell_6t
Xbit_r70_c226 bl_226 br_226 wl_70 vdd gnd cell_6t
Xbit_r71_c226 bl_226 br_226 wl_71 vdd gnd cell_6t
Xbit_r72_c226 bl_226 br_226 wl_72 vdd gnd cell_6t
Xbit_r73_c226 bl_226 br_226 wl_73 vdd gnd cell_6t
Xbit_r74_c226 bl_226 br_226 wl_74 vdd gnd cell_6t
Xbit_r75_c226 bl_226 br_226 wl_75 vdd gnd cell_6t
Xbit_r76_c226 bl_226 br_226 wl_76 vdd gnd cell_6t
Xbit_r77_c226 bl_226 br_226 wl_77 vdd gnd cell_6t
Xbit_r78_c226 bl_226 br_226 wl_78 vdd gnd cell_6t
Xbit_r79_c226 bl_226 br_226 wl_79 vdd gnd cell_6t
Xbit_r80_c226 bl_226 br_226 wl_80 vdd gnd cell_6t
Xbit_r81_c226 bl_226 br_226 wl_81 vdd gnd cell_6t
Xbit_r82_c226 bl_226 br_226 wl_82 vdd gnd cell_6t
Xbit_r83_c226 bl_226 br_226 wl_83 vdd gnd cell_6t
Xbit_r84_c226 bl_226 br_226 wl_84 vdd gnd cell_6t
Xbit_r85_c226 bl_226 br_226 wl_85 vdd gnd cell_6t
Xbit_r86_c226 bl_226 br_226 wl_86 vdd gnd cell_6t
Xbit_r87_c226 bl_226 br_226 wl_87 vdd gnd cell_6t
Xbit_r88_c226 bl_226 br_226 wl_88 vdd gnd cell_6t
Xbit_r89_c226 bl_226 br_226 wl_89 vdd gnd cell_6t
Xbit_r90_c226 bl_226 br_226 wl_90 vdd gnd cell_6t
Xbit_r91_c226 bl_226 br_226 wl_91 vdd gnd cell_6t
Xbit_r92_c226 bl_226 br_226 wl_92 vdd gnd cell_6t
Xbit_r93_c226 bl_226 br_226 wl_93 vdd gnd cell_6t
Xbit_r94_c226 bl_226 br_226 wl_94 vdd gnd cell_6t
Xbit_r95_c226 bl_226 br_226 wl_95 vdd gnd cell_6t
Xbit_r96_c226 bl_226 br_226 wl_96 vdd gnd cell_6t
Xbit_r97_c226 bl_226 br_226 wl_97 vdd gnd cell_6t
Xbit_r98_c226 bl_226 br_226 wl_98 vdd gnd cell_6t
Xbit_r99_c226 bl_226 br_226 wl_99 vdd gnd cell_6t
Xbit_r100_c226 bl_226 br_226 wl_100 vdd gnd cell_6t
Xbit_r101_c226 bl_226 br_226 wl_101 vdd gnd cell_6t
Xbit_r102_c226 bl_226 br_226 wl_102 vdd gnd cell_6t
Xbit_r103_c226 bl_226 br_226 wl_103 vdd gnd cell_6t
Xbit_r104_c226 bl_226 br_226 wl_104 vdd gnd cell_6t
Xbit_r105_c226 bl_226 br_226 wl_105 vdd gnd cell_6t
Xbit_r106_c226 bl_226 br_226 wl_106 vdd gnd cell_6t
Xbit_r107_c226 bl_226 br_226 wl_107 vdd gnd cell_6t
Xbit_r108_c226 bl_226 br_226 wl_108 vdd gnd cell_6t
Xbit_r109_c226 bl_226 br_226 wl_109 vdd gnd cell_6t
Xbit_r110_c226 bl_226 br_226 wl_110 vdd gnd cell_6t
Xbit_r111_c226 bl_226 br_226 wl_111 vdd gnd cell_6t
Xbit_r112_c226 bl_226 br_226 wl_112 vdd gnd cell_6t
Xbit_r113_c226 bl_226 br_226 wl_113 vdd gnd cell_6t
Xbit_r114_c226 bl_226 br_226 wl_114 vdd gnd cell_6t
Xbit_r115_c226 bl_226 br_226 wl_115 vdd gnd cell_6t
Xbit_r116_c226 bl_226 br_226 wl_116 vdd gnd cell_6t
Xbit_r117_c226 bl_226 br_226 wl_117 vdd gnd cell_6t
Xbit_r118_c226 bl_226 br_226 wl_118 vdd gnd cell_6t
Xbit_r119_c226 bl_226 br_226 wl_119 vdd gnd cell_6t
Xbit_r120_c226 bl_226 br_226 wl_120 vdd gnd cell_6t
Xbit_r121_c226 bl_226 br_226 wl_121 vdd gnd cell_6t
Xbit_r122_c226 bl_226 br_226 wl_122 vdd gnd cell_6t
Xbit_r123_c226 bl_226 br_226 wl_123 vdd gnd cell_6t
Xbit_r124_c226 bl_226 br_226 wl_124 vdd gnd cell_6t
Xbit_r125_c226 bl_226 br_226 wl_125 vdd gnd cell_6t
Xbit_r126_c226 bl_226 br_226 wl_126 vdd gnd cell_6t
Xbit_r127_c226 bl_226 br_226 wl_127 vdd gnd cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd cell_6t
Xbit_r1_c227 bl_227 br_227 wl_1 vdd gnd cell_6t
Xbit_r2_c227 bl_227 br_227 wl_2 vdd gnd cell_6t
Xbit_r3_c227 bl_227 br_227 wl_3 vdd gnd cell_6t
Xbit_r4_c227 bl_227 br_227 wl_4 vdd gnd cell_6t
Xbit_r5_c227 bl_227 br_227 wl_5 vdd gnd cell_6t
Xbit_r6_c227 bl_227 br_227 wl_6 vdd gnd cell_6t
Xbit_r7_c227 bl_227 br_227 wl_7 vdd gnd cell_6t
Xbit_r8_c227 bl_227 br_227 wl_8 vdd gnd cell_6t
Xbit_r9_c227 bl_227 br_227 wl_9 vdd gnd cell_6t
Xbit_r10_c227 bl_227 br_227 wl_10 vdd gnd cell_6t
Xbit_r11_c227 bl_227 br_227 wl_11 vdd gnd cell_6t
Xbit_r12_c227 bl_227 br_227 wl_12 vdd gnd cell_6t
Xbit_r13_c227 bl_227 br_227 wl_13 vdd gnd cell_6t
Xbit_r14_c227 bl_227 br_227 wl_14 vdd gnd cell_6t
Xbit_r15_c227 bl_227 br_227 wl_15 vdd gnd cell_6t
Xbit_r16_c227 bl_227 br_227 wl_16 vdd gnd cell_6t
Xbit_r17_c227 bl_227 br_227 wl_17 vdd gnd cell_6t
Xbit_r18_c227 bl_227 br_227 wl_18 vdd gnd cell_6t
Xbit_r19_c227 bl_227 br_227 wl_19 vdd gnd cell_6t
Xbit_r20_c227 bl_227 br_227 wl_20 vdd gnd cell_6t
Xbit_r21_c227 bl_227 br_227 wl_21 vdd gnd cell_6t
Xbit_r22_c227 bl_227 br_227 wl_22 vdd gnd cell_6t
Xbit_r23_c227 bl_227 br_227 wl_23 vdd gnd cell_6t
Xbit_r24_c227 bl_227 br_227 wl_24 vdd gnd cell_6t
Xbit_r25_c227 bl_227 br_227 wl_25 vdd gnd cell_6t
Xbit_r26_c227 bl_227 br_227 wl_26 vdd gnd cell_6t
Xbit_r27_c227 bl_227 br_227 wl_27 vdd gnd cell_6t
Xbit_r28_c227 bl_227 br_227 wl_28 vdd gnd cell_6t
Xbit_r29_c227 bl_227 br_227 wl_29 vdd gnd cell_6t
Xbit_r30_c227 bl_227 br_227 wl_30 vdd gnd cell_6t
Xbit_r31_c227 bl_227 br_227 wl_31 vdd gnd cell_6t
Xbit_r32_c227 bl_227 br_227 wl_32 vdd gnd cell_6t
Xbit_r33_c227 bl_227 br_227 wl_33 vdd gnd cell_6t
Xbit_r34_c227 bl_227 br_227 wl_34 vdd gnd cell_6t
Xbit_r35_c227 bl_227 br_227 wl_35 vdd gnd cell_6t
Xbit_r36_c227 bl_227 br_227 wl_36 vdd gnd cell_6t
Xbit_r37_c227 bl_227 br_227 wl_37 vdd gnd cell_6t
Xbit_r38_c227 bl_227 br_227 wl_38 vdd gnd cell_6t
Xbit_r39_c227 bl_227 br_227 wl_39 vdd gnd cell_6t
Xbit_r40_c227 bl_227 br_227 wl_40 vdd gnd cell_6t
Xbit_r41_c227 bl_227 br_227 wl_41 vdd gnd cell_6t
Xbit_r42_c227 bl_227 br_227 wl_42 vdd gnd cell_6t
Xbit_r43_c227 bl_227 br_227 wl_43 vdd gnd cell_6t
Xbit_r44_c227 bl_227 br_227 wl_44 vdd gnd cell_6t
Xbit_r45_c227 bl_227 br_227 wl_45 vdd gnd cell_6t
Xbit_r46_c227 bl_227 br_227 wl_46 vdd gnd cell_6t
Xbit_r47_c227 bl_227 br_227 wl_47 vdd gnd cell_6t
Xbit_r48_c227 bl_227 br_227 wl_48 vdd gnd cell_6t
Xbit_r49_c227 bl_227 br_227 wl_49 vdd gnd cell_6t
Xbit_r50_c227 bl_227 br_227 wl_50 vdd gnd cell_6t
Xbit_r51_c227 bl_227 br_227 wl_51 vdd gnd cell_6t
Xbit_r52_c227 bl_227 br_227 wl_52 vdd gnd cell_6t
Xbit_r53_c227 bl_227 br_227 wl_53 vdd gnd cell_6t
Xbit_r54_c227 bl_227 br_227 wl_54 vdd gnd cell_6t
Xbit_r55_c227 bl_227 br_227 wl_55 vdd gnd cell_6t
Xbit_r56_c227 bl_227 br_227 wl_56 vdd gnd cell_6t
Xbit_r57_c227 bl_227 br_227 wl_57 vdd gnd cell_6t
Xbit_r58_c227 bl_227 br_227 wl_58 vdd gnd cell_6t
Xbit_r59_c227 bl_227 br_227 wl_59 vdd gnd cell_6t
Xbit_r60_c227 bl_227 br_227 wl_60 vdd gnd cell_6t
Xbit_r61_c227 bl_227 br_227 wl_61 vdd gnd cell_6t
Xbit_r62_c227 bl_227 br_227 wl_62 vdd gnd cell_6t
Xbit_r63_c227 bl_227 br_227 wl_63 vdd gnd cell_6t
Xbit_r64_c227 bl_227 br_227 wl_64 vdd gnd cell_6t
Xbit_r65_c227 bl_227 br_227 wl_65 vdd gnd cell_6t
Xbit_r66_c227 bl_227 br_227 wl_66 vdd gnd cell_6t
Xbit_r67_c227 bl_227 br_227 wl_67 vdd gnd cell_6t
Xbit_r68_c227 bl_227 br_227 wl_68 vdd gnd cell_6t
Xbit_r69_c227 bl_227 br_227 wl_69 vdd gnd cell_6t
Xbit_r70_c227 bl_227 br_227 wl_70 vdd gnd cell_6t
Xbit_r71_c227 bl_227 br_227 wl_71 vdd gnd cell_6t
Xbit_r72_c227 bl_227 br_227 wl_72 vdd gnd cell_6t
Xbit_r73_c227 bl_227 br_227 wl_73 vdd gnd cell_6t
Xbit_r74_c227 bl_227 br_227 wl_74 vdd gnd cell_6t
Xbit_r75_c227 bl_227 br_227 wl_75 vdd gnd cell_6t
Xbit_r76_c227 bl_227 br_227 wl_76 vdd gnd cell_6t
Xbit_r77_c227 bl_227 br_227 wl_77 vdd gnd cell_6t
Xbit_r78_c227 bl_227 br_227 wl_78 vdd gnd cell_6t
Xbit_r79_c227 bl_227 br_227 wl_79 vdd gnd cell_6t
Xbit_r80_c227 bl_227 br_227 wl_80 vdd gnd cell_6t
Xbit_r81_c227 bl_227 br_227 wl_81 vdd gnd cell_6t
Xbit_r82_c227 bl_227 br_227 wl_82 vdd gnd cell_6t
Xbit_r83_c227 bl_227 br_227 wl_83 vdd gnd cell_6t
Xbit_r84_c227 bl_227 br_227 wl_84 vdd gnd cell_6t
Xbit_r85_c227 bl_227 br_227 wl_85 vdd gnd cell_6t
Xbit_r86_c227 bl_227 br_227 wl_86 vdd gnd cell_6t
Xbit_r87_c227 bl_227 br_227 wl_87 vdd gnd cell_6t
Xbit_r88_c227 bl_227 br_227 wl_88 vdd gnd cell_6t
Xbit_r89_c227 bl_227 br_227 wl_89 vdd gnd cell_6t
Xbit_r90_c227 bl_227 br_227 wl_90 vdd gnd cell_6t
Xbit_r91_c227 bl_227 br_227 wl_91 vdd gnd cell_6t
Xbit_r92_c227 bl_227 br_227 wl_92 vdd gnd cell_6t
Xbit_r93_c227 bl_227 br_227 wl_93 vdd gnd cell_6t
Xbit_r94_c227 bl_227 br_227 wl_94 vdd gnd cell_6t
Xbit_r95_c227 bl_227 br_227 wl_95 vdd gnd cell_6t
Xbit_r96_c227 bl_227 br_227 wl_96 vdd gnd cell_6t
Xbit_r97_c227 bl_227 br_227 wl_97 vdd gnd cell_6t
Xbit_r98_c227 bl_227 br_227 wl_98 vdd gnd cell_6t
Xbit_r99_c227 bl_227 br_227 wl_99 vdd gnd cell_6t
Xbit_r100_c227 bl_227 br_227 wl_100 vdd gnd cell_6t
Xbit_r101_c227 bl_227 br_227 wl_101 vdd gnd cell_6t
Xbit_r102_c227 bl_227 br_227 wl_102 vdd gnd cell_6t
Xbit_r103_c227 bl_227 br_227 wl_103 vdd gnd cell_6t
Xbit_r104_c227 bl_227 br_227 wl_104 vdd gnd cell_6t
Xbit_r105_c227 bl_227 br_227 wl_105 vdd gnd cell_6t
Xbit_r106_c227 bl_227 br_227 wl_106 vdd gnd cell_6t
Xbit_r107_c227 bl_227 br_227 wl_107 vdd gnd cell_6t
Xbit_r108_c227 bl_227 br_227 wl_108 vdd gnd cell_6t
Xbit_r109_c227 bl_227 br_227 wl_109 vdd gnd cell_6t
Xbit_r110_c227 bl_227 br_227 wl_110 vdd gnd cell_6t
Xbit_r111_c227 bl_227 br_227 wl_111 vdd gnd cell_6t
Xbit_r112_c227 bl_227 br_227 wl_112 vdd gnd cell_6t
Xbit_r113_c227 bl_227 br_227 wl_113 vdd gnd cell_6t
Xbit_r114_c227 bl_227 br_227 wl_114 vdd gnd cell_6t
Xbit_r115_c227 bl_227 br_227 wl_115 vdd gnd cell_6t
Xbit_r116_c227 bl_227 br_227 wl_116 vdd gnd cell_6t
Xbit_r117_c227 bl_227 br_227 wl_117 vdd gnd cell_6t
Xbit_r118_c227 bl_227 br_227 wl_118 vdd gnd cell_6t
Xbit_r119_c227 bl_227 br_227 wl_119 vdd gnd cell_6t
Xbit_r120_c227 bl_227 br_227 wl_120 vdd gnd cell_6t
Xbit_r121_c227 bl_227 br_227 wl_121 vdd gnd cell_6t
Xbit_r122_c227 bl_227 br_227 wl_122 vdd gnd cell_6t
Xbit_r123_c227 bl_227 br_227 wl_123 vdd gnd cell_6t
Xbit_r124_c227 bl_227 br_227 wl_124 vdd gnd cell_6t
Xbit_r125_c227 bl_227 br_227 wl_125 vdd gnd cell_6t
Xbit_r126_c227 bl_227 br_227 wl_126 vdd gnd cell_6t
Xbit_r127_c227 bl_227 br_227 wl_127 vdd gnd cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd cell_6t
Xbit_r1_c228 bl_228 br_228 wl_1 vdd gnd cell_6t
Xbit_r2_c228 bl_228 br_228 wl_2 vdd gnd cell_6t
Xbit_r3_c228 bl_228 br_228 wl_3 vdd gnd cell_6t
Xbit_r4_c228 bl_228 br_228 wl_4 vdd gnd cell_6t
Xbit_r5_c228 bl_228 br_228 wl_5 vdd gnd cell_6t
Xbit_r6_c228 bl_228 br_228 wl_6 vdd gnd cell_6t
Xbit_r7_c228 bl_228 br_228 wl_7 vdd gnd cell_6t
Xbit_r8_c228 bl_228 br_228 wl_8 vdd gnd cell_6t
Xbit_r9_c228 bl_228 br_228 wl_9 vdd gnd cell_6t
Xbit_r10_c228 bl_228 br_228 wl_10 vdd gnd cell_6t
Xbit_r11_c228 bl_228 br_228 wl_11 vdd gnd cell_6t
Xbit_r12_c228 bl_228 br_228 wl_12 vdd gnd cell_6t
Xbit_r13_c228 bl_228 br_228 wl_13 vdd gnd cell_6t
Xbit_r14_c228 bl_228 br_228 wl_14 vdd gnd cell_6t
Xbit_r15_c228 bl_228 br_228 wl_15 vdd gnd cell_6t
Xbit_r16_c228 bl_228 br_228 wl_16 vdd gnd cell_6t
Xbit_r17_c228 bl_228 br_228 wl_17 vdd gnd cell_6t
Xbit_r18_c228 bl_228 br_228 wl_18 vdd gnd cell_6t
Xbit_r19_c228 bl_228 br_228 wl_19 vdd gnd cell_6t
Xbit_r20_c228 bl_228 br_228 wl_20 vdd gnd cell_6t
Xbit_r21_c228 bl_228 br_228 wl_21 vdd gnd cell_6t
Xbit_r22_c228 bl_228 br_228 wl_22 vdd gnd cell_6t
Xbit_r23_c228 bl_228 br_228 wl_23 vdd gnd cell_6t
Xbit_r24_c228 bl_228 br_228 wl_24 vdd gnd cell_6t
Xbit_r25_c228 bl_228 br_228 wl_25 vdd gnd cell_6t
Xbit_r26_c228 bl_228 br_228 wl_26 vdd gnd cell_6t
Xbit_r27_c228 bl_228 br_228 wl_27 vdd gnd cell_6t
Xbit_r28_c228 bl_228 br_228 wl_28 vdd gnd cell_6t
Xbit_r29_c228 bl_228 br_228 wl_29 vdd gnd cell_6t
Xbit_r30_c228 bl_228 br_228 wl_30 vdd gnd cell_6t
Xbit_r31_c228 bl_228 br_228 wl_31 vdd gnd cell_6t
Xbit_r32_c228 bl_228 br_228 wl_32 vdd gnd cell_6t
Xbit_r33_c228 bl_228 br_228 wl_33 vdd gnd cell_6t
Xbit_r34_c228 bl_228 br_228 wl_34 vdd gnd cell_6t
Xbit_r35_c228 bl_228 br_228 wl_35 vdd gnd cell_6t
Xbit_r36_c228 bl_228 br_228 wl_36 vdd gnd cell_6t
Xbit_r37_c228 bl_228 br_228 wl_37 vdd gnd cell_6t
Xbit_r38_c228 bl_228 br_228 wl_38 vdd gnd cell_6t
Xbit_r39_c228 bl_228 br_228 wl_39 vdd gnd cell_6t
Xbit_r40_c228 bl_228 br_228 wl_40 vdd gnd cell_6t
Xbit_r41_c228 bl_228 br_228 wl_41 vdd gnd cell_6t
Xbit_r42_c228 bl_228 br_228 wl_42 vdd gnd cell_6t
Xbit_r43_c228 bl_228 br_228 wl_43 vdd gnd cell_6t
Xbit_r44_c228 bl_228 br_228 wl_44 vdd gnd cell_6t
Xbit_r45_c228 bl_228 br_228 wl_45 vdd gnd cell_6t
Xbit_r46_c228 bl_228 br_228 wl_46 vdd gnd cell_6t
Xbit_r47_c228 bl_228 br_228 wl_47 vdd gnd cell_6t
Xbit_r48_c228 bl_228 br_228 wl_48 vdd gnd cell_6t
Xbit_r49_c228 bl_228 br_228 wl_49 vdd gnd cell_6t
Xbit_r50_c228 bl_228 br_228 wl_50 vdd gnd cell_6t
Xbit_r51_c228 bl_228 br_228 wl_51 vdd gnd cell_6t
Xbit_r52_c228 bl_228 br_228 wl_52 vdd gnd cell_6t
Xbit_r53_c228 bl_228 br_228 wl_53 vdd gnd cell_6t
Xbit_r54_c228 bl_228 br_228 wl_54 vdd gnd cell_6t
Xbit_r55_c228 bl_228 br_228 wl_55 vdd gnd cell_6t
Xbit_r56_c228 bl_228 br_228 wl_56 vdd gnd cell_6t
Xbit_r57_c228 bl_228 br_228 wl_57 vdd gnd cell_6t
Xbit_r58_c228 bl_228 br_228 wl_58 vdd gnd cell_6t
Xbit_r59_c228 bl_228 br_228 wl_59 vdd gnd cell_6t
Xbit_r60_c228 bl_228 br_228 wl_60 vdd gnd cell_6t
Xbit_r61_c228 bl_228 br_228 wl_61 vdd gnd cell_6t
Xbit_r62_c228 bl_228 br_228 wl_62 vdd gnd cell_6t
Xbit_r63_c228 bl_228 br_228 wl_63 vdd gnd cell_6t
Xbit_r64_c228 bl_228 br_228 wl_64 vdd gnd cell_6t
Xbit_r65_c228 bl_228 br_228 wl_65 vdd gnd cell_6t
Xbit_r66_c228 bl_228 br_228 wl_66 vdd gnd cell_6t
Xbit_r67_c228 bl_228 br_228 wl_67 vdd gnd cell_6t
Xbit_r68_c228 bl_228 br_228 wl_68 vdd gnd cell_6t
Xbit_r69_c228 bl_228 br_228 wl_69 vdd gnd cell_6t
Xbit_r70_c228 bl_228 br_228 wl_70 vdd gnd cell_6t
Xbit_r71_c228 bl_228 br_228 wl_71 vdd gnd cell_6t
Xbit_r72_c228 bl_228 br_228 wl_72 vdd gnd cell_6t
Xbit_r73_c228 bl_228 br_228 wl_73 vdd gnd cell_6t
Xbit_r74_c228 bl_228 br_228 wl_74 vdd gnd cell_6t
Xbit_r75_c228 bl_228 br_228 wl_75 vdd gnd cell_6t
Xbit_r76_c228 bl_228 br_228 wl_76 vdd gnd cell_6t
Xbit_r77_c228 bl_228 br_228 wl_77 vdd gnd cell_6t
Xbit_r78_c228 bl_228 br_228 wl_78 vdd gnd cell_6t
Xbit_r79_c228 bl_228 br_228 wl_79 vdd gnd cell_6t
Xbit_r80_c228 bl_228 br_228 wl_80 vdd gnd cell_6t
Xbit_r81_c228 bl_228 br_228 wl_81 vdd gnd cell_6t
Xbit_r82_c228 bl_228 br_228 wl_82 vdd gnd cell_6t
Xbit_r83_c228 bl_228 br_228 wl_83 vdd gnd cell_6t
Xbit_r84_c228 bl_228 br_228 wl_84 vdd gnd cell_6t
Xbit_r85_c228 bl_228 br_228 wl_85 vdd gnd cell_6t
Xbit_r86_c228 bl_228 br_228 wl_86 vdd gnd cell_6t
Xbit_r87_c228 bl_228 br_228 wl_87 vdd gnd cell_6t
Xbit_r88_c228 bl_228 br_228 wl_88 vdd gnd cell_6t
Xbit_r89_c228 bl_228 br_228 wl_89 vdd gnd cell_6t
Xbit_r90_c228 bl_228 br_228 wl_90 vdd gnd cell_6t
Xbit_r91_c228 bl_228 br_228 wl_91 vdd gnd cell_6t
Xbit_r92_c228 bl_228 br_228 wl_92 vdd gnd cell_6t
Xbit_r93_c228 bl_228 br_228 wl_93 vdd gnd cell_6t
Xbit_r94_c228 bl_228 br_228 wl_94 vdd gnd cell_6t
Xbit_r95_c228 bl_228 br_228 wl_95 vdd gnd cell_6t
Xbit_r96_c228 bl_228 br_228 wl_96 vdd gnd cell_6t
Xbit_r97_c228 bl_228 br_228 wl_97 vdd gnd cell_6t
Xbit_r98_c228 bl_228 br_228 wl_98 vdd gnd cell_6t
Xbit_r99_c228 bl_228 br_228 wl_99 vdd gnd cell_6t
Xbit_r100_c228 bl_228 br_228 wl_100 vdd gnd cell_6t
Xbit_r101_c228 bl_228 br_228 wl_101 vdd gnd cell_6t
Xbit_r102_c228 bl_228 br_228 wl_102 vdd gnd cell_6t
Xbit_r103_c228 bl_228 br_228 wl_103 vdd gnd cell_6t
Xbit_r104_c228 bl_228 br_228 wl_104 vdd gnd cell_6t
Xbit_r105_c228 bl_228 br_228 wl_105 vdd gnd cell_6t
Xbit_r106_c228 bl_228 br_228 wl_106 vdd gnd cell_6t
Xbit_r107_c228 bl_228 br_228 wl_107 vdd gnd cell_6t
Xbit_r108_c228 bl_228 br_228 wl_108 vdd gnd cell_6t
Xbit_r109_c228 bl_228 br_228 wl_109 vdd gnd cell_6t
Xbit_r110_c228 bl_228 br_228 wl_110 vdd gnd cell_6t
Xbit_r111_c228 bl_228 br_228 wl_111 vdd gnd cell_6t
Xbit_r112_c228 bl_228 br_228 wl_112 vdd gnd cell_6t
Xbit_r113_c228 bl_228 br_228 wl_113 vdd gnd cell_6t
Xbit_r114_c228 bl_228 br_228 wl_114 vdd gnd cell_6t
Xbit_r115_c228 bl_228 br_228 wl_115 vdd gnd cell_6t
Xbit_r116_c228 bl_228 br_228 wl_116 vdd gnd cell_6t
Xbit_r117_c228 bl_228 br_228 wl_117 vdd gnd cell_6t
Xbit_r118_c228 bl_228 br_228 wl_118 vdd gnd cell_6t
Xbit_r119_c228 bl_228 br_228 wl_119 vdd gnd cell_6t
Xbit_r120_c228 bl_228 br_228 wl_120 vdd gnd cell_6t
Xbit_r121_c228 bl_228 br_228 wl_121 vdd gnd cell_6t
Xbit_r122_c228 bl_228 br_228 wl_122 vdd gnd cell_6t
Xbit_r123_c228 bl_228 br_228 wl_123 vdd gnd cell_6t
Xbit_r124_c228 bl_228 br_228 wl_124 vdd gnd cell_6t
Xbit_r125_c228 bl_228 br_228 wl_125 vdd gnd cell_6t
Xbit_r126_c228 bl_228 br_228 wl_126 vdd gnd cell_6t
Xbit_r127_c228 bl_228 br_228 wl_127 vdd gnd cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd cell_6t
Xbit_r1_c229 bl_229 br_229 wl_1 vdd gnd cell_6t
Xbit_r2_c229 bl_229 br_229 wl_2 vdd gnd cell_6t
Xbit_r3_c229 bl_229 br_229 wl_3 vdd gnd cell_6t
Xbit_r4_c229 bl_229 br_229 wl_4 vdd gnd cell_6t
Xbit_r5_c229 bl_229 br_229 wl_5 vdd gnd cell_6t
Xbit_r6_c229 bl_229 br_229 wl_6 vdd gnd cell_6t
Xbit_r7_c229 bl_229 br_229 wl_7 vdd gnd cell_6t
Xbit_r8_c229 bl_229 br_229 wl_8 vdd gnd cell_6t
Xbit_r9_c229 bl_229 br_229 wl_9 vdd gnd cell_6t
Xbit_r10_c229 bl_229 br_229 wl_10 vdd gnd cell_6t
Xbit_r11_c229 bl_229 br_229 wl_11 vdd gnd cell_6t
Xbit_r12_c229 bl_229 br_229 wl_12 vdd gnd cell_6t
Xbit_r13_c229 bl_229 br_229 wl_13 vdd gnd cell_6t
Xbit_r14_c229 bl_229 br_229 wl_14 vdd gnd cell_6t
Xbit_r15_c229 bl_229 br_229 wl_15 vdd gnd cell_6t
Xbit_r16_c229 bl_229 br_229 wl_16 vdd gnd cell_6t
Xbit_r17_c229 bl_229 br_229 wl_17 vdd gnd cell_6t
Xbit_r18_c229 bl_229 br_229 wl_18 vdd gnd cell_6t
Xbit_r19_c229 bl_229 br_229 wl_19 vdd gnd cell_6t
Xbit_r20_c229 bl_229 br_229 wl_20 vdd gnd cell_6t
Xbit_r21_c229 bl_229 br_229 wl_21 vdd gnd cell_6t
Xbit_r22_c229 bl_229 br_229 wl_22 vdd gnd cell_6t
Xbit_r23_c229 bl_229 br_229 wl_23 vdd gnd cell_6t
Xbit_r24_c229 bl_229 br_229 wl_24 vdd gnd cell_6t
Xbit_r25_c229 bl_229 br_229 wl_25 vdd gnd cell_6t
Xbit_r26_c229 bl_229 br_229 wl_26 vdd gnd cell_6t
Xbit_r27_c229 bl_229 br_229 wl_27 vdd gnd cell_6t
Xbit_r28_c229 bl_229 br_229 wl_28 vdd gnd cell_6t
Xbit_r29_c229 bl_229 br_229 wl_29 vdd gnd cell_6t
Xbit_r30_c229 bl_229 br_229 wl_30 vdd gnd cell_6t
Xbit_r31_c229 bl_229 br_229 wl_31 vdd gnd cell_6t
Xbit_r32_c229 bl_229 br_229 wl_32 vdd gnd cell_6t
Xbit_r33_c229 bl_229 br_229 wl_33 vdd gnd cell_6t
Xbit_r34_c229 bl_229 br_229 wl_34 vdd gnd cell_6t
Xbit_r35_c229 bl_229 br_229 wl_35 vdd gnd cell_6t
Xbit_r36_c229 bl_229 br_229 wl_36 vdd gnd cell_6t
Xbit_r37_c229 bl_229 br_229 wl_37 vdd gnd cell_6t
Xbit_r38_c229 bl_229 br_229 wl_38 vdd gnd cell_6t
Xbit_r39_c229 bl_229 br_229 wl_39 vdd gnd cell_6t
Xbit_r40_c229 bl_229 br_229 wl_40 vdd gnd cell_6t
Xbit_r41_c229 bl_229 br_229 wl_41 vdd gnd cell_6t
Xbit_r42_c229 bl_229 br_229 wl_42 vdd gnd cell_6t
Xbit_r43_c229 bl_229 br_229 wl_43 vdd gnd cell_6t
Xbit_r44_c229 bl_229 br_229 wl_44 vdd gnd cell_6t
Xbit_r45_c229 bl_229 br_229 wl_45 vdd gnd cell_6t
Xbit_r46_c229 bl_229 br_229 wl_46 vdd gnd cell_6t
Xbit_r47_c229 bl_229 br_229 wl_47 vdd gnd cell_6t
Xbit_r48_c229 bl_229 br_229 wl_48 vdd gnd cell_6t
Xbit_r49_c229 bl_229 br_229 wl_49 vdd gnd cell_6t
Xbit_r50_c229 bl_229 br_229 wl_50 vdd gnd cell_6t
Xbit_r51_c229 bl_229 br_229 wl_51 vdd gnd cell_6t
Xbit_r52_c229 bl_229 br_229 wl_52 vdd gnd cell_6t
Xbit_r53_c229 bl_229 br_229 wl_53 vdd gnd cell_6t
Xbit_r54_c229 bl_229 br_229 wl_54 vdd gnd cell_6t
Xbit_r55_c229 bl_229 br_229 wl_55 vdd gnd cell_6t
Xbit_r56_c229 bl_229 br_229 wl_56 vdd gnd cell_6t
Xbit_r57_c229 bl_229 br_229 wl_57 vdd gnd cell_6t
Xbit_r58_c229 bl_229 br_229 wl_58 vdd gnd cell_6t
Xbit_r59_c229 bl_229 br_229 wl_59 vdd gnd cell_6t
Xbit_r60_c229 bl_229 br_229 wl_60 vdd gnd cell_6t
Xbit_r61_c229 bl_229 br_229 wl_61 vdd gnd cell_6t
Xbit_r62_c229 bl_229 br_229 wl_62 vdd gnd cell_6t
Xbit_r63_c229 bl_229 br_229 wl_63 vdd gnd cell_6t
Xbit_r64_c229 bl_229 br_229 wl_64 vdd gnd cell_6t
Xbit_r65_c229 bl_229 br_229 wl_65 vdd gnd cell_6t
Xbit_r66_c229 bl_229 br_229 wl_66 vdd gnd cell_6t
Xbit_r67_c229 bl_229 br_229 wl_67 vdd gnd cell_6t
Xbit_r68_c229 bl_229 br_229 wl_68 vdd gnd cell_6t
Xbit_r69_c229 bl_229 br_229 wl_69 vdd gnd cell_6t
Xbit_r70_c229 bl_229 br_229 wl_70 vdd gnd cell_6t
Xbit_r71_c229 bl_229 br_229 wl_71 vdd gnd cell_6t
Xbit_r72_c229 bl_229 br_229 wl_72 vdd gnd cell_6t
Xbit_r73_c229 bl_229 br_229 wl_73 vdd gnd cell_6t
Xbit_r74_c229 bl_229 br_229 wl_74 vdd gnd cell_6t
Xbit_r75_c229 bl_229 br_229 wl_75 vdd gnd cell_6t
Xbit_r76_c229 bl_229 br_229 wl_76 vdd gnd cell_6t
Xbit_r77_c229 bl_229 br_229 wl_77 vdd gnd cell_6t
Xbit_r78_c229 bl_229 br_229 wl_78 vdd gnd cell_6t
Xbit_r79_c229 bl_229 br_229 wl_79 vdd gnd cell_6t
Xbit_r80_c229 bl_229 br_229 wl_80 vdd gnd cell_6t
Xbit_r81_c229 bl_229 br_229 wl_81 vdd gnd cell_6t
Xbit_r82_c229 bl_229 br_229 wl_82 vdd gnd cell_6t
Xbit_r83_c229 bl_229 br_229 wl_83 vdd gnd cell_6t
Xbit_r84_c229 bl_229 br_229 wl_84 vdd gnd cell_6t
Xbit_r85_c229 bl_229 br_229 wl_85 vdd gnd cell_6t
Xbit_r86_c229 bl_229 br_229 wl_86 vdd gnd cell_6t
Xbit_r87_c229 bl_229 br_229 wl_87 vdd gnd cell_6t
Xbit_r88_c229 bl_229 br_229 wl_88 vdd gnd cell_6t
Xbit_r89_c229 bl_229 br_229 wl_89 vdd gnd cell_6t
Xbit_r90_c229 bl_229 br_229 wl_90 vdd gnd cell_6t
Xbit_r91_c229 bl_229 br_229 wl_91 vdd gnd cell_6t
Xbit_r92_c229 bl_229 br_229 wl_92 vdd gnd cell_6t
Xbit_r93_c229 bl_229 br_229 wl_93 vdd gnd cell_6t
Xbit_r94_c229 bl_229 br_229 wl_94 vdd gnd cell_6t
Xbit_r95_c229 bl_229 br_229 wl_95 vdd gnd cell_6t
Xbit_r96_c229 bl_229 br_229 wl_96 vdd gnd cell_6t
Xbit_r97_c229 bl_229 br_229 wl_97 vdd gnd cell_6t
Xbit_r98_c229 bl_229 br_229 wl_98 vdd gnd cell_6t
Xbit_r99_c229 bl_229 br_229 wl_99 vdd gnd cell_6t
Xbit_r100_c229 bl_229 br_229 wl_100 vdd gnd cell_6t
Xbit_r101_c229 bl_229 br_229 wl_101 vdd gnd cell_6t
Xbit_r102_c229 bl_229 br_229 wl_102 vdd gnd cell_6t
Xbit_r103_c229 bl_229 br_229 wl_103 vdd gnd cell_6t
Xbit_r104_c229 bl_229 br_229 wl_104 vdd gnd cell_6t
Xbit_r105_c229 bl_229 br_229 wl_105 vdd gnd cell_6t
Xbit_r106_c229 bl_229 br_229 wl_106 vdd gnd cell_6t
Xbit_r107_c229 bl_229 br_229 wl_107 vdd gnd cell_6t
Xbit_r108_c229 bl_229 br_229 wl_108 vdd gnd cell_6t
Xbit_r109_c229 bl_229 br_229 wl_109 vdd gnd cell_6t
Xbit_r110_c229 bl_229 br_229 wl_110 vdd gnd cell_6t
Xbit_r111_c229 bl_229 br_229 wl_111 vdd gnd cell_6t
Xbit_r112_c229 bl_229 br_229 wl_112 vdd gnd cell_6t
Xbit_r113_c229 bl_229 br_229 wl_113 vdd gnd cell_6t
Xbit_r114_c229 bl_229 br_229 wl_114 vdd gnd cell_6t
Xbit_r115_c229 bl_229 br_229 wl_115 vdd gnd cell_6t
Xbit_r116_c229 bl_229 br_229 wl_116 vdd gnd cell_6t
Xbit_r117_c229 bl_229 br_229 wl_117 vdd gnd cell_6t
Xbit_r118_c229 bl_229 br_229 wl_118 vdd gnd cell_6t
Xbit_r119_c229 bl_229 br_229 wl_119 vdd gnd cell_6t
Xbit_r120_c229 bl_229 br_229 wl_120 vdd gnd cell_6t
Xbit_r121_c229 bl_229 br_229 wl_121 vdd gnd cell_6t
Xbit_r122_c229 bl_229 br_229 wl_122 vdd gnd cell_6t
Xbit_r123_c229 bl_229 br_229 wl_123 vdd gnd cell_6t
Xbit_r124_c229 bl_229 br_229 wl_124 vdd gnd cell_6t
Xbit_r125_c229 bl_229 br_229 wl_125 vdd gnd cell_6t
Xbit_r126_c229 bl_229 br_229 wl_126 vdd gnd cell_6t
Xbit_r127_c229 bl_229 br_229 wl_127 vdd gnd cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd cell_6t
Xbit_r1_c230 bl_230 br_230 wl_1 vdd gnd cell_6t
Xbit_r2_c230 bl_230 br_230 wl_2 vdd gnd cell_6t
Xbit_r3_c230 bl_230 br_230 wl_3 vdd gnd cell_6t
Xbit_r4_c230 bl_230 br_230 wl_4 vdd gnd cell_6t
Xbit_r5_c230 bl_230 br_230 wl_5 vdd gnd cell_6t
Xbit_r6_c230 bl_230 br_230 wl_6 vdd gnd cell_6t
Xbit_r7_c230 bl_230 br_230 wl_7 vdd gnd cell_6t
Xbit_r8_c230 bl_230 br_230 wl_8 vdd gnd cell_6t
Xbit_r9_c230 bl_230 br_230 wl_9 vdd gnd cell_6t
Xbit_r10_c230 bl_230 br_230 wl_10 vdd gnd cell_6t
Xbit_r11_c230 bl_230 br_230 wl_11 vdd gnd cell_6t
Xbit_r12_c230 bl_230 br_230 wl_12 vdd gnd cell_6t
Xbit_r13_c230 bl_230 br_230 wl_13 vdd gnd cell_6t
Xbit_r14_c230 bl_230 br_230 wl_14 vdd gnd cell_6t
Xbit_r15_c230 bl_230 br_230 wl_15 vdd gnd cell_6t
Xbit_r16_c230 bl_230 br_230 wl_16 vdd gnd cell_6t
Xbit_r17_c230 bl_230 br_230 wl_17 vdd gnd cell_6t
Xbit_r18_c230 bl_230 br_230 wl_18 vdd gnd cell_6t
Xbit_r19_c230 bl_230 br_230 wl_19 vdd gnd cell_6t
Xbit_r20_c230 bl_230 br_230 wl_20 vdd gnd cell_6t
Xbit_r21_c230 bl_230 br_230 wl_21 vdd gnd cell_6t
Xbit_r22_c230 bl_230 br_230 wl_22 vdd gnd cell_6t
Xbit_r23_c230 bl_230 br_230 wl_23 vdd gnd cell_6t
Xbit_r24_c230 bl_230 br_230 wl_24 vdd gnd cell_6t
Xbit_r25_c230 bl_230 br_230 wl_25 vdd gnd cell_6t
Xbit_r26_c230 bl_230 br_230 wl_26 vdd gnd cell_6t
Xbit_r27_c230 bl_230 br_230 wl_27 vdd gnd cell_6t
Xbit_r28_c230 bl_230 br_230 wl_28 vdd gnd cell_6t
Xbit_r29_c230 bl_230 br_230 wl_29 vdd gnd cell_6t
Xbit_r30_c230 bl_230 br_230 wl_30 vdd gnd cell_6t
Xbit_r31_c230 bl_230 br_230 wl_31 vdd gnd cell_6t
Xbit_r32_c230 bl_230 br_230 wl_32 vdd gnd cell_6t
Xbit_r33_c230 bl_230 br_230 wl_33 vdd gnd cell_6t
Xbit_r34_c230 bl_230 br_230 wl_34 vdd gnd cell_6t
Xbit_r35_c230 bl_230 br_230 wl_35 vdd gnd cell_6t
Xbit_r36_c230 bl_230 br_230 wl_36 vdd gnd cell_6t
Xbit_r37_c230 bl_230 br_230 wl_37 vdd gnd cell_6t
Xbit_r38_c230 bl_230 br_230 wl_38 vdd gnd cell_6t
Xbit_r39_c230 bl_230 br_230 wl_39 vdd gnd cell_6t
Xbit_r40_c230 bl_230 br_230 wl_40 vdd gnd cell_6t
Xbit_r41_c230 bl_230 br_230 wl_41 vdd gnd cell_6t
Xbit_r42_c230 bl_230 br_230 wl_42 vdd gnd cell_6t
Xbit_r43_c230 bl_230 br_230 wl_43 vdd gnd cell_6t
Xbit_r44_c230 bl_230 br_230 wl_44 vdd gnd cell_6t
Xbit_r45_c230 bl_230 br_230 wl_45 vdd gnd cell_6t
Xbit_r46_c230 bl_230 br_230 wl_46 vdd gnd cell_6t
Xbit_r47_c230 bl_230 br_230 wl_47 vdd gnd cell_6t
Xbit_r48_c230 bl_230 br_230 wl_48 vdd gnd cell_6t
Xbit_r49_c230 bl_230 br_230 wl_49 vdd gnd cell_6t
Xbit_r50_c230 bl_230 br_230 wl_50 vdd gnd cell_6t
Xbit_r51_c230 bl_230 br_230 wl_51 vdd gnd cell_6t
Xbit_r52_c230 bl_230 br_230 wl_52 vdd gnd cell_6t
Xbit_r53_c230 bl_230 br_230 wl_53 vdd gnd cell_6t
Xbit_r54_c230 bl_230 br_230 wl_54 vdd gnd cell_6t
Xbit_r55_c230 bl_230 br_230 wl_55 vdd gnd cell_6t
Xbit_r56_c230 bl_230 br_230 wl_56 vdd gnd cell_6t
Xbit_r57_c230 bl_230 br_230 wl_57 vdd gnd cell_6t
Xbit_r58_c230 bl_230 br_230 wl_58 vdd gnd cell_6t
Xbit_r59_c230 bl_230 br_230 wl_59 vdd gnd cell_6t
Xbit_r60_c230 bl_230 br_230 wl_60 vdd gnd cell_6t
Xbit_r61_c230 bl_230 br_230 wl_61 vdd gnd cell_6t
Xbit_r62_c230 bl_230 br_230 wl_62 vdd gnd cell_6t
Xbit_r63_c230 bl_230 br_230 wl_63 vdd gnd cell_6t
Xbit_r64_c230 bl_230 br_230 wl_64 vdd gnd cell_6t
Xbit_r65_c230 bl_230 br_230 wl_65 vdd gnd cell_6t
Xbit_r66_c230 bl_230 br_230 wl_66 vdd gnd cell_6t
Xbit_r67_c230 bl_230 br_230 wl_67 vdd gnd cell_6t
Xbit_r68_c230 bl_230 br_230 wl_68 vdd gnd cell_6t
Xbit_r69_c230 bl_230 br_230 wl_69 vdd gnd cell_6t
Xbit_r70_c230 bl_230 br_230 wl_70 vdd gnd cell_6t
Xbit_r71_c230 bl_230 br_230 wl_71 vdd gnd cell_6t
Xbit_r72_c230 bl_230 br_230 wl_72 vdd gnd cell_6t
Xbit_r73_c230 bl_230 br_230 wl_73 vdd gnd cell_6t
Xbit_r74_c230 bl_230 br_230 wl_74 vdd gnd cell_6t
Xbit_r75_c230 bl_230 br_230 wl_75 vdd gnd cell_6t
Xbit_r76_c230 bl_230 br_230 wl_76 vdd gnd cell_6t
Xbit_r77_c230 bl_230 br_230 wl_77 vdd gnd cell_6t
Xbit_r78_c230 bl_230 br_230 wl_78 vdd gnd cell_6t
Xbit_r79_c230 bl_230 br_230 wl_79 vdd gnd cell_6t
Xbit_r80_c230 bl_230 br_230 wl_80 vdd gnd cell_6t
Xbit_r81_c230 bl_230 br_230 wl_81 vdd gnd cell_6t
Xbit_r82_c230 bl_230 br_230 wl_82 vdd gnd cell_6t
Xbit_r83_c230 bl_230 br_230 wl_83 vdd gnd cell_6t
Xbit_r84_c230 bl_230 br_230 wl_84 vdd gnd cell_6t
Xbit_r85_c230 bl_230 br_230 wl_85 vdd gnd cell_6t
Xbit_r86_c230 bl_230 br_230 wl_86 vdd gnd cell_6t
Xbit_r87_c230 bl_230 br_230 wl_87 vdd gnd cell_6t
Xbit_r88_c230 bl_230 br_230 wl_88 vdd gnd cell_6t
Xbit_r89_c230 bl_230 br_230 wl_89 vdd gnd cell_6t
Xbit_r90_c230 bl_230 br_230 wl_90 vdd gnd cell_6t
Xbit_r91_c230 bl_230 br_230 wl_91 vdd gnd cell_6t
Xbit_r92_c230 bl_230 br_230 wl_92 vdd gnd cell_6t
Xbit_r93_c230 bl_230 br_230 wl_93 vdd gnd cell_6t
Xbit_r94_c230 bl_230 br_230 wl_94 vdd gnd cell_6t
Xbit_r95_c230 bl_230 br_230 wl_95 vdd gnd cell_6t
Xbit_r96_c230 bl_230 br_230 wl_96 vdd gnd cell_6t
Xbit_r97_c230 bl_230 br_230 wl_97 vdd gnd cell_6t
Xbit_r98_c230 bl_230 br_230 wl_98 vdd gnd cell_6t
Xbit_r99_c230 bl_230 br_230 wl_99 vdd gnd cell_6t
Xbit_r100_c230 bl_230 br_230 wl_100 vdd gnd cell_6t
Xbit_r101_c230 bl_230 br_230 wl_101 vdd gnd cell_6t
Xbit_r102_c230 bl_230 br_230 wl_102 vdd gnd cell_6t
Xbit_r103_c230 bl_230 br_230 wl_103 vdd gnd cell_6t
Xbit_r104_c230 bl_230 br_230 wl_104 vdd gnd cell_6t
Xbit_r105_c230 bl_230 br_230 wl_105 vdd gnd cell_6t
Xbit_r106_c230 bl_230 br_230 wl_106 vdd gnd cell_6t
Xbit_r107_c230 bl_230 br_230 wl_107 vdd gnd cell_6t
Xbit_r108_c230 bl_230 br_230 wl_108 vdd gnd cell_6t
Xbit_r109_c230 bl_230 br_230 wl_109 vdd gnd cell_6t
Xbit_r110_c230 bl_230 br_230 wl_110 vdd gnd cell_6t
Xbit_r111_c230 bl_230 br_230 wl_111 vdd gnd cell_6t
Xbit_r112_c230 bl_230 br_230 wl_112 vdd gnd cell_6t
Xbit_r113_c230 bl_230 br_230 wl_113 vdd gnd cell_6t
Xbit_r114_c230 bl_230 br_230 wl_114 vdd gnd cell_6t
Xbit_r115_c230 bl_230 br_230 wl_115 vdd gnd cell_6t
Xbit_r116_c230 bl_230 br_230 wl_116 vdd gnd cell_6t
Xbit_r117_c230 bl_230 br_230 wl_117 vdd gnd cell_6t
Xbit_r118_c230 bl_230 br_230 wl_118 vdd gnd cell_6t
Xbit_r119_c230 bl_230 br_230 wl_119 vdd gnd cell_6t
Xbit_r120_c230 bl_230 br_230 wl_120 vdd gnd cell_6t
Xbit_r121_c230 bl_230 br_230 wl_121 vdd gnd cell_6t
Xbit_r122_c230 bl_230 br_230 wl_122 vdd gnd cell_6t
Xbit_r123_c230 bl_230 br_230 wl_123 vdd gnd cell_6t
Xbit_r124_c230 bl_230 br_230 wl_124 vdd gnd cell_6t
Xbit_r125_c230 bl_230 br_230 wl_125 vdd gnd cell_6t
Xbit_r126_c230 bl_230 br_230 wl_126 vdd gnd cell_6t
Xbit_r127_c230 bl_230 br_230 wl_127 vdd gnd cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd cell_6t
Xbit_r1_c231 bl_231 br_231 wl_1 vdd gnd cell_6t
Xbit_r2_c231 bl_231 br_231 wl_2 vdd gnd cell_6t
Xbit_r3_c231 bl_231 br_231 wl_3 vdd gnd cell_6t
Xbit_r4_c231 bl_231 br_231 wl_4 vdd gnd cell_6t
Xbit_r5_c231 bl_231 br_231 wl_5 vdd gnd cell_6t
Xbit_r6_c231 bl_231 br_231 wl_6 vdd gnd cell_6t
Xbit_r7_c231 bl_231 br_231 wl_7 vdd gnd cell_6t
Xbit_r8_c231 bl_231 br_231 wl_8 vdd gnd cell_6t
Xbit_r9_c231 bl_231 br_231 wl_9 vdd gnd cell_6t
Xbit_r10_c231 bl_231 br_231 wl_10 vdd gnd cell_6t
Xbit_r11_c231 bl_231 br_231 wl_11 vdd gnd cell_6t
Xbit_r12_c231 bl_231 br_231 wl_12 vdd gnd cell_6t
Xbit_r13_c231 bl_231 br_231 wl_13 vdd gnd cell_6t
Xbit_r14_c231 bl_231 br_231 wl_14 vdd gnd cell_6t
Xbit_r15_c231 bl_231 br_231 wl_15 vdd gnd cell_6t
Xbit_r16_c231 bl_231 br_231 wl_16 vdd gnd cell_6t
Xbit_r17_c231 bl_231 br_231 wl_17 vdd gnd cell_6t
Xbit_r18_c231 bl_231 br_231 wl_18 vdd gnd cell_6t
Xbit_r19_c231 bl_231 br_231 wl_19 vdd gnd cell_6t
Xbit_r20_c231 bl_231 br_231 wl_20 vdd gnd cell_6t
Xbit_r21_c231 bl_231 br_231 wl_21 vdd gnd cell_6t
Xbit_r22_c231 bl_231 br_231 wl_22 vdd gnd cell_6t
Xbit_r23_c231 bl_231 br_231 wl_23 vdd gnd cell_6t
Xbit_r24_c231 bl_231 br_231 wl_24 vdd gnd cell_6t
Xbit_r25_c231 bl_231 br_231 wl_25 vdd gnd cell_6t
Xbit_r26_c231 bl_231 br_231 wl_26 vdd gnd cell_6t
Xbit_r27_c231 bl_231 br_231 wl_27 vdd gnd cell_6t
Xbit_r28_c231 bl_231 br_231 wl_28 vdd gnd cell_6t
Xbit_r29_c231 bl_231 br_231 wl_29 vdd gnd cell_6t
Xbit_r30_c231 bl_231 br_231 wl_30 vdd gnd cell_6t
Xbit_r31_c231 bl_231 br_231 wl_31 vdd gnd cell_6t
Xbit_r32_c231 bl_231 br_231 wl_32 vdd gnd cell_6t
Xbit_r33_c231 bl_231 br_231 wl_33 vdd gnd cell_6t
Xbit_r34_c231 bl_231 br_231 wl_34 vdd gnd cell_6t
Xbit_r35_c231 bl_231 br_231 wl_35 vdd gnd cell_6t
Xbit_r36_c231 bl_231 br_231 wl_36 vdd gnd cell_6t
Xbit_r37_c231 bl_231 br_231 wl_37 vdd gnd cell_6t
Xbit_r38_c231 bl_231 br_231 wl_38 vdd gnd cell_6t
Xbit_r39_c231 bl_231 br_231 wl_39 vdd gnd cell_6t
Xbit_r40_c231 bl_231 br_231 wl_40 vdd gnd cell_6t
Xbit_r41_c231 bl_231 br_231 wl_41 vdd gnd cell_6t
Xbit_r42_c231 bl_231 br_231 wl_42 vdd gnd cell_6t
Xbit_r43_c231 bl_231 br_231 wl_43 vdd gnd cell_6t
Xbit_r44_c231 bl_231 br_231 wl_44 vdd gnd cell_6t
Xbit_r45_c231 bl_231 br_231 wl_45 vdd gnd cell_6t
Xbit_r46_c231 bl_231 br_231 wl_46 vdd gnd cell_6t
Xbit_r47_c231 bl_231 br_231 wl_47 vdd gnd cell_6t
Xbit_r48_c231 bl_231 br_231 wl_48 vdd gnd cell_6t
Xbit_r49_c231 bl_231 br_231 wl_49 vdd gnd cell_6t
Xbit_r50_c231 bl_231 br_231 wl_50 vdd gnd cell_6t
Xbit_r51_c231 bl_231 br_231 wl_51 vdd gnd cell_6t
Xbit_r52_c231 bl_231 br_231 wl_52 vdd gnd cell_6t
Xbit_r53_c231 bl_231 br_231 wl_53 vdd gnd cell_6t
Xbit_r54_c231 bl_231 br_231 wl_54 vdd gnd cell_6t
Xbit_r55_c231 bl_231 br_231 wl_55 vdd gnd cell_6t
Xbit_r56_c231 bl_231 br_231 wl_56 vdd gnd cell_6t
Xbit_r57_c231 bl_231 br_231 wl_57 vdd gnd cell_6t
Xbit_r58_c231 bl_231 br_231 wl_58 vdd gnd cell_6t
Xbit_r59_c231 bl_231 br_231 wl_59 vdd gnd cell_6t
Xbit_r60_c231 bl_231 br_231 wl_60 vdd gnd cell_6t
Xbit_r61_c231 bl_231 br_231 wl_61 vdd gnd cell_6t
Xbit_r62_c231 bl_231 br_231 wl_62 vdd gnd cell_6t
Xbit_r63_c231 bl_231 br_231 wl_63 vdd gnd cell_6t
Xbit_r64_c231 bl_231 br_231 wl_64 vdd gnd cell_6t
Xbit_r65_c231 bl_231 br_231 wl_65 vdd gnd cell_6t
Xbit_r66_c231 bl_231 br_231 wl_66 vdd gnd cell_6t
Xbit_r67_c231 bl_231 br_231 wl_67 vdd gnd cell_6t
Xbit_r68_c231 bl_231 br_231 wl_68 vdd gnd cell_6t
Xbit_r69_c231 bl_231 br_231 wl_69 vdd gnd cell_6t
Xbit_r70_c231 bl_231 br_231 wl_70 vdd gnd cell_6t
Xbit_r71_c231 bl_231 br_231 wl_71 vdd gnd cell_6t
Xbit_r72_c231 bl_231 br_231 wl_72 vdd gnd cell_6t
Xbit_r73_c231 bl_231 br_231 wl_73 vdd gnd cell_6t
Xbit_r74_c231 bl_231 br_231 wl_74 vdd gnd cell_6t
Xbit_r75_c231 bl_231 br_231 wl_75 vdd gnd cell_6t
Xbit_r76_c231 bl_231 br_231 wl_76 vdd gnd cell_6t
Xbit_r77_c231 bl_231 br_231 wl_77 vdd gnd cell_6t
Xbit_r78_c231 bl_231 br_231 wl_78 vdd gnd cell_6t
Xbit_r79_c231 bl_231 br_231 wl_79 vdd gnd cell_6t
Xbit_r80_c231 bl_231 br_231 wl_80 vdd gnd cell_6t
Xbit_r81_c231 bl_231 br_231 wl_81 vdd gnd cell_6t
Xbit_r82_c231 bl_231 br_231 wl_82 vdd gnd cell_6t
Xbit_r83_c231 bl_231 br_231 wl_83 vdd gnd cell_6t
Xbit_r84_c231 bl_231 br_231 wl_84 vdd gnd cell_6t
Xbit_r85_c231 bl_231 br_231 wl_85 vdd gnd cell_6t
Xbit_r86_c231 bl_231 br_231 wl_86 vdd gnd cell_6t
Xbit_r87_c231 bl_231 br_231 wl_87 vdd gnd cell_6t
Xbit_r88_c231 bl_231 br_231 wl_88 vdd gnd cell_6t
Xbit_r89_c231 bl_231 br_231 wl_89 vdd gnd cell_6t
Xbit_r90_c231 bl_231 br_231 wl_90 vdd gnd cell_6t
Xbit_r91_c231 bl_231 br_231 wl_91 vdd gnd cell_6t
Xbit_r92_c231 bl_231 br_231 wl_92 vdd gnd cell_6t
Xbit_r93_c231 bl_231 br_231 wl_93 vdd gnd cell_6t
Xbit_r94_c231 bl_231 br_231 wl_94 vdd gnd cell_6t
Xbit_r95_c231 bl_231 br_231 wl_95 vdd gnd cell_6t
Xbit_r96_c231 bl_231 br_231 wl_96 vdd gnd cell_6t
Xbit_r97_c231 bl_231 br_231 wl_97 vdd gnd cell_6t
Xbit_r98_c231 bl_231 br_231 wl_98 vdd gnd cell_6t
Xbit_r99_c231 bl_231 br_231 wl_99 vdd gnd cell_6t
Xbit_r100_c231 bl_231 br_231 wl_100 vdd gnd cell_6t
Xbit_r101_c231 bl_231 br_231 wl_101 vdd gnd cell_6t
Xbit_r102_c231 bl_231 br_231 wl_102 vdd gnd cell_6t
Xbit_r103_c231 bl_231 br_231 wl_103 vdd gnd cell_6t
Xbit_r104_c231 bl_231 br_231 wl_104 vdd gnd cell_6t
Xbit_r105_c231 bl_231 br_231 wl_105 vdd gnd cell_6t
Xbit_r106_c231 bl_231 br_231 wl_106 vdd gnd cell_6t
Xbit_r107_c231 bl_231 br_231 wl_107 vdd gnd cell_6t
Xbit_r108_c231 bl_231 br_231 wl_108 vdd gnd cell_6t
Xbit_r109_c231 bl_231 br_231 wl_109 vdd gnd cell_6t
Xbit_r110_c231 bl_231 br_231 wl_110 vdd gnd cell_6t
Xbit_r111_c231 bl_231 br_231 wl_111 vdd gnd cell_6t
Xbit_r112_c231 bl_231 br_231 wl_112 vdd gnd cell_6t
Xbit_r113_c231 bl_231 br_231 wl_113 vdd gnd cell_6t
Xbit_r114_c231 bl_231 br_231 wl_114 vdd gnd cell_6t
Xbit_r115_c231 bl_231 br_231 wl_115 vdd gnd cell_6t
Xbit_r116_c231 bl_231 br_231 wl_116 vdd gnd cell_6t
Xbit_r117_c231 bl_231 br_231 wl_117 vdd gnd cell_6t
Xbit_r118_c231 bl_231 br_231 wl_118 vdd gnd cell_6t
Xbit_r119_c231 bl_231 br_231 wl_119 vdd gnd cell_6t
Xbit_r120_c231 bl_231 br_231 wl_120 vdd gnd cell_6t
Xbit_r121_c231 bl_231 br_231 wl_121 vdd gnd cell_6t
Xbit_r122_c231 bl_231 br_231 wl_122 vdd gnd cell_6t
Xbit_r123_c231 bl_231 br_231 wl_123 vdd gnd cell_6t
Xbit_r124_c231 bl_231 br_231 wl_124 vdd gnd cell_6t
Xbit_r125_c231 bl_231 br_231 wl_125 vdd gnd cell_6t
Xbit_r126_c231 bl_231 br_231 wl_126 vdd gnd cell_6t
Xbit_r127_c231 bl_231 br_231 wl_127 vdd gnd cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd cell_6t
Xbit_r1_c232 bl_232 br_232 wl_1 vdd gnd cell_6t
Xbit_r2_c232 bl_232 br_232 wl_2 vdd gnd cell_6t
Xbit_r3_c232 bl_232 br_232 wl_3 vdd gnd cell_6t
Xbit_r4_c232 bl_232 br_232 wl_4 vdd gnd cell_6t
Xbit_r5_c232 bl_232 br_232 wl_5 vdd gnd cell_6t
Xbit_r6_c232 bl_232 br_232 wl_6 vdd gnd cell_6t
Xbit_r7_c232 bl_232 br_232 wl_7 vdd gnd cell_6t
Xbit_r8_c232 bl_232 br_232 wl_8 vdd gnd cell_6t
Xbit_r9_c232 bl_232 br_232 wl_9 vdd gnd cell_6t
Xbit_r10_c232 bl_232 br_232 wl_10 vdd gnd cell_6t
Xbit_r11_c232 bl_232 br_232 wl_11 vdd gnd cell_6t
Xbit_r12_c232 bl_232 br_232 wl_12 vdd gnd cell_6t
Xbit_r13_c232 bl_232 br_232 wl_13 vdd gnd cell_6t
Xbit_r14_c232 bl_232 br_232 wl_14 vdd gnd cell_6t
Xbit_r15_c232 bl_232 br_232 wl_15 vdd gnd cell_6t
Xbit_r16_c232 bl_232 br_232 wl_16 vdd gnd cell_6t
Xbit_r17_c232 bl_232 br_232 wl_17 vdd gnd cell_6t
Xbit_r18_c232 bl_232 br_232 wl_18 vdd gnd cell_6t
Xbit_r19_c232 bl_232 br_232 wl_19 vdd gnd cell_6t
Xbit_r20_c232 bl_232 br_232 wl_20 vdd gnd cell_6t
Xbit_r21_c232 bl_232 br_232 wl_21 vdd gnd cell_6t
Xbit_r22_c232 bl_232 br_232 wl_22 vdd gnd cell_6t
Xbit_r23_c232 bl_232 br_232 wl_23 vdd gnd cell_6t
Xbit_r24_c232 bl_232 br_232 wl_24 vdd gnd cell_6t
Xbit_r25_c232 bl_232 br_232 wl_25 vdd gnd cell_6t
Xbit_r26_c232 bl_232 br_232 wl_26 vdd gnd cell_6t
Xbit_r27_c232 bl_232 br_232 wl_27 vdd gnd cell_6t
Xbit_r28_c232 bl_232 br_232 wl_28 vdd gnd cell_6t
Xbit_r29_c232 bl_232 br_232 wl_29 vdd gnd cell_6t
Xbit_r30_c232 bl_232 br_232 wl_30 vdd gnd cell_6t
Xbit_r31_c232 bl_232 br_232 wl_31 vdd gnd cell_6t
Xbit_r32_c232 bl_232 br_232 wl_32 vdd gnd cell_6t
Xbit_r33_c232 bl_232 br_232 wl_33 vdd gnd cell_6t
Xbit_r34_c232 bl_232 br_232 wl_34 vdd gnd cell_6t
Xbit_r35_c232 bl_232 br_232 wl_35 vdd gnd cell_6t
Xbit_r36_c232 bl_232 br_232 wl_36 vdd gnd cell_6t
Xbit_r37_c232 bl_232 br_232 wl_37 vdd gnd cell_6t
Xbit_r38_c232 bl_232 br_232 wl_38 vdd gnd cell_6t
Xbit_r39_c232 bl_232 br_232 wl_39 vdd gnd cell_6t
Xbit_r40_c232 bl_232 br_232 wl_40 vdd gnd cell_6t
Xbit_r41_c232 bl_232 br_232 wl_41 vdd gnd cell_6t
Xbit_r42_c232 bl_232 br_232 wl_42 vdd gnd cell_6t
Xbit_r43_c232 bl_232 br_232 wl_43 vdd gnd cell_6t
Xbit_r44_c232 bl_232 br_232 wl_44 vdd gnd cell_6t
Xbit_r45_c232 bl_232 br_232 wl_45 vdd gnd cell_6t
Xbit_r46_c232 bl_232 br_232 wl_46 vdd gnd cell_6t
Xbit_r47_c232 bl_232 br_232 wl_47 vdd gnd cell_6t
Xbit_r48_c232 bl_232 br_232 wl_48 vdd gnd cell_6t
Xbit_r49_c232 bl_232 br_232 wl_49 vdd gnd cell_6t
Xbit_r50_c232 bl_232 br_232 wl_50 vdd gnd cell_6t
Xbit_r51_c232 bl_232 br_232 wl_51 vdd gnd cell_6t
Xbit_r52_c232 bl_232 br_232 wl_52 vdd gnd cell_6t
Xbit_r53_c232 bl_232 br_232 wl_53 vdd gnd cell_6t
Xbit_r54_c232 bl_232 br_232 wl_54 vdd gnd cell_6t
Xbit_r55_c232 bl_232 br_232 wl_55 vdd gnd cell_6t
Xbit_r56_c232 bl_232 br_232 wl_56 vdd gnd cell_6t
Xbit_r57_c232 bl_232 br_232 wl_57 vdd gnd cell_6t
Xbit_r58_c232 bl_232 br_232 wl_58 vdd gnd cell_6t
Xbit_r59_c232 bl_232 br_232 wl_59 vdd gnd cell_6t
Xbit_r60_c232 bl_232 br_232 wl_60 vdd gnd cell_6t
Xbit_r61_c232 bl_232 br_232 wl_61 vdd gnd cell_6t
Xbit_r62_c232 bl_232 br_232 wl_62 vdd gnd cell_6t
Xbit_r63_c232 bl_232 br_232 wl_63 vdd gnd cell_6t
Xbit_r64_c232 bl_232 br_232 wl_64 vdd gnd cell_6t
Xbit_r65_c232 bl_232 br_232 wl_65 vdd gnd cell_6t
Xbit_r66_c232 bl_232 br_232 wl_66 vdd gnd cell_6t
Xbit_r67_c232 bl_232 br_232 wl_67 vdd gnd cell_6t
Xbit_r68_c232 bl_232 br_232 wl_68 vdd gnd cell_6t
Xbit_r69_c232 bl_232 br_232 wl_69 vdd gnd cell_6t
Xbit_r70_c232 bl_232 br_232 wl_70 vdd gnd cell_6t
Xbit_r71_c232 bl_232 br_232 wl_71 vdd gnd cell_6t
Xbit_r72_c232 bl_232 br_232 wl_72 vdd gnd cell_6t
Xbit_r73_c232 bl_232 br_232 wl_73 vdd gnd cell_6t
Xbit_r74_c232 bl_232 br_232 wl_74 vdd gnd cell_6t
Xbit_r75_c232 bl_232 br_232 wl_75 vdd gnd cell_6t
Xbit_r76_c232 bl_232 br_232 wl_76 vdd gnd cell_6t
Xbit_r77_c232 bl_232 br_232 wl_77 vdd gnd cell_6t
Xbit_r78_c232 bl_232 br_232 wl_78 vdd gnd cell_6t
Xbit_r79_c232 bl_232 br_232 wl_79 vdd gnd cell_6t
Xbit_r80_c232 bl_232 br_232 wl_80 vdd gnd cell_6t
Xbit_r81_c232 bl_232 br_232 wl_81 vdd gnd cell_6t
Xbit_r82_c232 bl_232 br_232 wl_82 vdd gnd cell_6t
Xbit_r83_c232 bl_232 br_232 wl_83 vdd gnd cell_6t
Xbit_r84_c232 bl_232 br_232 wl_84 vdd gnd cell_6t
Xbit_r85_c232 bl_232 br_232 wl_85 vdd gnd cell_6t
Xbit_r86_c232 bl_232 br_232 wl_86 vdd gnd cell_6t
Xbit_r87_c232 bl_232 br_232 wl_87 vdd gnd cell_6t
Xbit_r88_c232 bl_232 br_232 wl_88 vdd gnd cell_6t
Xbit_r89_c232 bl_232 br_232 wl_89 vdd gnd cell_6t
Xbit_r90_c232 bl_232 br_232 wl_90 vdd gnd cell_6t
Xbit_r91_c232 bl_232 br_232 wl_91 vdd gnd cell_6t
Xbit_r92_c232 bl_232 br_232 wl_92 vdd gnd cell_6t
Xbit_r93_c232 bl_232 br_232 wl_93 vdd gnd cell_6t
Xbit_r94_c232 bl_232 br_232 wl_94 vdd gnd cell_6t
Xbit_r95_c232 bl_232 br_232 wl_95 vdd gnd cell_6t
Xbit_r96_c232 bl_232 br_232 wl_96 vdd gnd cell_6t
Xbit_r97_c232 bl_232 br_232 wl_97 vdd gnd cell_6t
Xbit_r98_c232 bl_232 br_232 wl_98 vdd gnd cell_6t
Xbit_r99_c232 bl_232 br_232 wl_99 vdd gnd cell_6t
Xbit_r100_c232 bl_232 br_232 wl_100 vdd gnd cell_6t
Xbit_r101_c232 bl_232 br_232 wl_101 vdd gnd cell_6t
Xbit_r102_c232 bl_232 br_232 wl_102 vdd gnd cell_6t
Xbit_r103_c232 bl_232 br_232 wl_103 vdd gnd cell_6t
Xbit_r104_c232 bl_232 br_232 wl_104 vdd gnd cell_6t
Xbit_r105_c232 bl_232 br_232 wl_105 vdd gnd cell_6t
Xbit_r106_c232 bl_232 br_232 wl_106 vdd gnd cell_6t
Xbit_r107_c232 bl_232 br_232 wl_107 vdd gnd cell_6t
Xbit_r108_c232 bl_232 br_232 wl_108 vdd gnd cell_6t
Xbit_r109_c232 bl_232 br_232 wl_109 vdd gnd cell_6t
Xbit_r110_c232 bl_232 br_232 wl_110 vdd gnd cell_6t
Xbit_r111_c232 bl_232 br_232 wl_111 vdd gnd cell_6t
Xbit_r112_c232 bl_232 br_232 wl_112 vdd gnd cell_6t
Xbit_r113_c232 bl_232 br_232 wl_113 vdd gnd cell_6t
Xbit_r114_c232 bl_232 br_232 wl_114 vdd gnd cell_6t
Xbit_r115_c232 bl_232 br_232 wl_115 vdd gnd cell_6t
Xbit_r116_c232 bl_232 br_232 wl_116 vdd gnd cell_6t
Xbit_r117_c232 bl_232 br_232 wl_117 vdd gnd cell_6t
Xbit_r118_c232 bl_232 br_232 wl_118 vdd gnd cell_6t
Xbit_r119_c232 bl_232 br_232 wl_119 vdd gnd cell_6t
Xbit_r120_c232 bl_232 br_232 wl_120 vdd gnd cell_6t
Xbit_r121_c232 bl_232 br_232 wl_121 vdd gnd cell_6t
Xbit_r122_c232 bl_232 br_232 wl_122 vdd gnd cell_6t
Xbit_r123_c232 bl_232 br_232 wl_123 vdd gnd cell_6t
Xbit_r124_c232 bl_232 br_232 wl_124 vdd gnd cell_6t
Xbit_r125_c232 bl_232 br_232 wl_125 vdd gnd cell_6t
Xbit_r126_c232 bl_232 br_232 wl_126 vdd gnd cell_6t
Xbit_r127_c232 bl_232 br_232 wl_127 vdd gnd cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd cell_6t
Xbit_r1_c233 bl_233 br_233 wl_1 vdd gnd cell_6t
Xbit_r2_c233 bl_233 br_233 wl_2 vdd gnd cell_6t
Xbit_r3_c233 bl_233 br_233 wl_3 vdd gnd cell_6t
Xbit_r4_c233 bl_233 br_233 wl_4 vdd gnd cell_6t
Xbit_r5_c233 bl_233 br_233 wl_5 vdd gnd cell_6t
Xbit_r6_c233 bl_233 br_233 wl_6 vdd gnd cell_6t
Xbit_r7_c233 bl_233 br_233 wl_7 vdd gnd cell_6t
Xbit_r8_c233 bl_233 br_233 wl_8 vdd gnd cell_6t
Xbit_r9_c233 bl_233 br_233 wl_9 vdd gnd cell_6t
Xbit_r10_c233 bl_233 br_233 wl_10 vdd gnd cell_6t
Xbit_r11_c233 bl_233 br_233 wl_11 vdd gnd cell_6t
Xbit_r12_c233 bl_233 br_233 wl_12 vdd gnd cell_6t
Xbit_r13_c233 bl_233 br_233 wl_13 vdd gnd cell_6t
Xbit_r14_c233 bl_233 br_233 wl_14 vdd gnd cell_6t
Xbit_r15_c233 bl_233 br_233 wl_15 vdd gnd cell_6t
Xbit_r16_c233 bl_233 br_233 wl_16 vdd gnd cell_6t
Xbit_r17_c233 bl_233 br_233 wl_17 vdd gnd cell_6t
Xbit_r18_c233 bl_233 br_233 wl_18 vdd gnd cell_6t
Xbit_r19_c233 bl_233 br_233 wl_19 vdd gnd cell_6t
Xbit_r20_c233 bl_233 br_233 wl_20 vdd gnd cell_6t
Xbit_r21_c233 bl_233 br_233 wl_21 vdd gnd cell_6t
Xbit_r22_c233 bl_233 br_233 wl_22 vdd gnd cell_6t
Xbit_r23_c233 bl_233 br_233 wl_23 vdd gnd cell_6t
Xbit_r24_c233 bl_233 br_233 wl_24 vdd gnd cell_6t
Xbit_r25_c233 bl_233 br_233 wl_25 vdd gnd cell_6t
Xbit_r26_c233 bl_233 br_233 wl_26 vdd gnd cell_6t
Xbit_r27_c233 bl_233 br_233 wl_27 vdd gnd cell_6t
Xbit_r28_c233 bl_233 br_233 wl_28 vdd gnd cell_6t
Xbit_r29_c233 bl_233 br_233 wl_29 vdd gnd cell_6t
Xbit_r30_c233 bl_233 br_233 wl_30 vdd gnd cell_6t
Xbit_r31_c233 bl_233 br_233 wl_31 vdd gnd cell_6t
Xbit_r32_c233 bl_233 br_233 wl_32 vdd gnd cell_6t
Xbit_r33_c233 bl_233 br_233 wl_33 vdd gnd cell_6t
Xbit_r34_c233 bl_233 br_233 wl_34 vdd gnd cell_6t
Xbit_r35_c233 bl_233 br_233 wl_35 vdd gnd cell_6t
Xbit_r36_c233 bl_233 br_233 wl_36 vdd gnd cell_6t
Xbit_r37_c233 bl_233 br_233 wl_37 vdd gnd cell_6t
Xbit_r38_c233 bl_233 br_233 wl_38 vdd gnd cell_6t
Xbit_r39_c233 bl_233 br_233 wl_39 vdd gnd cell_6t
Xbit_r40_c233 bl_233 br_233 wl_40 vdd gnd cell_6t
Xbit_r41_c233 bl_233 br_233 wl_41 vdd gnd cell_6t
Xbit_r42_c233 bl_233 br_233 wl_42 vdd gnd cell_6t
Xbit_r43_c233 bl_233 br_233 wl_43 vdd gnd cell_6t
Xbit_r44_c233 bl_233 br_233 wl_44 vdd gnd cell_6t
Xbit_r45_c233 bl_233 br_233 wl_45 vdd gnd cell_6t
Xbit_r46_c233 bl_233 br_233 wl_46 vdd gnd cell_6t
Xbit_r47_c233 bl_233 br_233 wl_47 vdd gnd cell_6t
Xbit_r48_c233 bl_233 br_233 wl_48 vdd gnd cell_6t
Xbit_r49_c233 bl_233 br_233 wl_49 vdd gnd cell_6t
Xbit_r50_c233 bl_233 br_233 wl_50 vdd gnd cell_6t
Xbit_r51_c233 bl_233 br_233 wl_51 vdd gnd cell_6t
Xbit_r52_c233 bl_233 br_233 wl_52 vdd gnd cell_6t
Xbit_r53_c233 bl_233 br_233 wl_53 vdd gnd cell_6t
Xbit_r54_c233 bl_233 br_233 wl_54 vdd gnd cell_6t
Xbit_r55_c233 bl_233 br_233 wl_55 vdd gnd cell_6t
Xbit_r56_c233 bl_233 br_233 wl_56 vdd gnd cell_6t
Xbit_r57_c233 bl_233 br_233 wl_57 vdd gnd cell_6t
Xbit_r58_c233 bl_233 br_233 wl_58 vdd gnd cell_6t
Xbit_r59_c233 bl_233 br_233 wl_59 vdd gnd cell_6t
Xbit_r60_c233 bl_233 br_233 wl_60 vdd gnd cell_6t
Xbit_r61_c233 bl_233 br_233 wl_61 vdd gnd cell_6t
Xbit_r62_c233 bl_233 br_233 wl_62 vdd gnd cell_6t
Xbit_r63_c233 bl_233 br_233 wl_63 vdd gnd cell_6t
Xbit_r64_c233 bl_233 br_233 wl_64 vdd gnd cell_6t
Xbit_r65_c233 bl_233 br_233 wl_65 vdd gnd cell_6t
Xbit_r66_c233 bl_233 br_233 wl_66 vdd gnd cell_6t
Xbit_r67_c233 bl_233 br_233 wl_67 vdd gnd cell_6t
Xbit_r68_c233 bl_233 br_233 wl_68 vdd gnd cell_6t
Xbit_r69_c233 bl_233 br_233 wl_69 vdd gnd cell_6t
Xbit_r70_c233 bl_233 br_233 wl_70 vdd gnd cell_6t
Xbit_r71_c233 bl_233 br_233 wl_71 vdd gnd cell_6t
Xbit_r72_c233 bl_233 br_233 wl_72 vdd gnd cell_6t
Xbit_r73_c233 bl_233 br_233 wl_73 vdd gnd cell_6t
Xbit_r74_c233 bl_233 br_233 wl_74 vdd gnd cell_6t
Xbit_r75_c233 bl_233 br_233 wl_75 vdd gnd cell_6t
Xbit_r76_c233 bl_233 br_233 wl_76 vdd gnd cell_6t
Xbit_r77_c233 bl_233 br_233 wl_77 vdd gnd cell_6t
Xbit_r78_c233 bl_233 br_233 wl_78 vdd gnd cell_6t
Xbit_r79_c233 bl_233 br_233 wl_79 vdd gnd cell_6t
Xbit_r80_c233 bl_233 br_233 wl_80 vdd gnd cell_6t
Xbit_r81_c233 bl_233 br_233 wl_81 vdd gnd cell_6t
Xbit_r82_c233 bl_233 br_233 wl_82 vdd gnd cell_6t
Xbit_r83_c233 bl_233 br_233 wl_83 vdd gnd cell_6t
Xbit_r84_c233 bl_233 br_233 wl_84 vdd gnd cell_6t
Xbit_r85_c233 bl_233 br_233 wl_85 vdd gnd cell_6t
Xbit_r86_c233 bl_233 br_233 wl_86 vdd gnd cell_6t
Xbit_r87_c233 bl_233 br_233 wl_87 vdd gnd cell_6t
Xbit_r88_c233 bl_233 br_233 wl_88 vdd gnd cell_6t
Xbit_r89_c233 bl_233 br_233 wl_89 vdd gnd cell_6t
Xbit_r90_c233 bl_233 br_233 wl_90 vdd gnd cell_6t
Xbit_r91_c233 bl_233 br_233 wl_91 vdd gnd cell_6t
Xbit_r92_c233 bl_233 br_233 wl_92 vdd gnd cell_6t
Xbit_r93_c233 bl_233 br_233 wl_93 vdd gnd cell_6t
Xbit_r94_c233 bl_233 br_233 wl_94 vdd gnd cell_6t
Xbit_r95_c233 bl_233 br_233 wl_95 vdd gnd cell_6t
Xbit_r96_c233 bl_233 br_233 wl_96 vdd gnd cell_6t
Xbit_r97_c233 bl_233 br_233 wl_97 vdd gnd cell_6t
Xbit_r98_c233 bl_233 br_233 wl_98 vdd gnd cell_6t
Xbit_r99_c233 bl_233 br_233 wl_99 vdd gnd cell_6t
Xbit_r100_c233 bl_233 br_233 wl_100 vdd gnd cell_6t
Xbit_r101_c233 bl_233 br_233 wl_101 vdd gnd cell_6t
Xbit_r102_c233 bl_233 br_233 wl_102 vdd gnd cell_6t
Xbit_r103_c233 bl_233 br_233 wl_103 vdd gnd cell_6t
Xbit_r104_c233 bl_233 br_233 wl_104 vdd gnd cell_6t
Xbit_r105_c233 bl_233 br_233 wl_105 vdd gnd cell_6t
Xbit_r106_c233 bl_233 br_233 wl_106 vdd gnd cell_6t
Xbit_r107_c233 bl_233 br_233 wl_107 vdd gnd cell_6t
Xbit_r108_c233 bl_233 br_233 wl_108 vdd gnd cell_6t
Xbit_r109_c233 bl_233 br_233 wl_109 vdd gnd cell_6t
Xbit_r110_c233 bl_233 br_233 wl_110 vdd gnd cell_6t
Xbit_r111_c233 bl_233 br_233 wl_111 vdd gnd cell_6t
Xbit_r112_c233 bl_233 br_233 wl_112 vdd gnd cell_6t
Xbit_r113_c233 bl_233 br_233 wl_113 vdd gnd cell_6t
Xbit_r114_c233 bl_233 br_233 wl_114 vdd gnd cell_6t
Xbit_r115_c233 bl_233 br_233 wl_115 vdd gnd cell_6t
Xbit_r116_c233 bl_233 br_233 wl_116 vdd gnd cell_6t
Xbit_r117_c233 bl_233 br_233 wl_117 vdd gnd cell_6t
Xbit_r118_c233 bl_233 br_233 wl_118 vdd gnd cell_6t
Xbit_r119_c233 bl_233 br_233 wl_119 vdd gnd cell_6t
Xbit_r120_c233 bl_233 br_233 wl_120 vdd gnd cell_6t
Xbit_r121_c233 bl_233 br_233 wl_121 vdd gnd cell_6t
Xbit_r122_c233 bl_233 br_233 wl_122 vdd gnd cell_6t
Xbit_r123_c233 bl_233 br_233 wl_123 vdd gnd cell_6t
Xbit_r124_c233 bl_233 br_233 wl_124 vdd gnd cell_6t
Xbit_r125_c233 bl_233 br_233 wl_125 vdd gnd cell_6t
Xbit_r126_c233 bl_233 br_233 wl_126 vdd gnd cell_6t
Xbit_r127_c233 bl_233 br_233 wl_127 vdd gnd cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd cell_6t
Xbit_r1_c234 bl_234 br_234 wl_1 vdd gnd cell_6t
Xbit_r2_c234 bl_234 br_234 wl_2 vdd gnd cell_6t
Xbit_r3_c234 bl_234 br_234 wl_3 vdd gnd cell_6t
Xbit_r4_c234 bl_234 br_234 wl_4 vdd gnd cell_6t
Xbit_r5_c234 bl_234 br_234 wl_5 vdd gnd cell_6t
Xbit_r6_c234 bl_234 br_234 wl_6 vdd gnd cell_6t
Xbit_r7_c234 bl_234 br_234 wl_7 vdd gnd cell_6t
Xbit_r8_c234 bl_234 br_234 wl_8 vdd gnd cell_6t
Xbit_r9_c234 bl_234 br_234 wl_9 vdd gnd cell_6t
Xbit_r10_c234 bl_234 br_234 wl_10 vdd gnd cell_6t
Xbit_r11_c234 bl_234 br_234 wl_11 vdd gnd cell_6t
Xbit_r12_c234 bl_234 br_234 wl_12 vdd gnd cell_6t
Xbit_r13_c234 bl_234 br_234 wl_13 vdd gnd cell_6t
Xbit_r14_c234 bl_234 br_234 wl_14 vdd gnd cell_6t
Xbit_r15_c234 bl_234 br_234 wl_15 vdd gnd cell_6t
Xbit_r16_c234 bl_234 br_234 wl_16 vdd gnd cell_6t
Xbit_r17_c234 bl_234 br_234 wl_17 vdd gnd cell_6t
Xbit_r18_c234 bl_234 br_234 wl_18 vdd gnd cell_6t
Xbit_r19_c234 bl_234 br_234 wl_19 vdd gnd cell_6t
Xbit_r20_c234 bl_234 br_234 wl_20 vdd gnd cell_6t
Xbit_r21_c234 bl_234 br_234 wl_21 vdd gnd cell_6t
Xbit_r22_c234 bl_234 br_234 wl_22 vdd gnd cell_6t
Xbit_r23_c234 bl_234 br_234 wl_23 vdd gnd cell_6t
Xbit_r24_c234 bl_234 br_234 wl_24 vdd gnd cell_6t
Xbit_r25_c234 bl_234 br_234 wl_25 vdd gnd cell_6t
Xbit_r26_c234 bl_234 br_234 wl_26 vdd gnd cell_6t
Xbit_r27_c234 bl_234 br_234 wl_27 vdd gnd cell_6t
Xbit_r28_c234 bl_234 br_234 wl_28 vdd gnd cell_6t
Xbit_r29_c234 bl_234 br_234 wl_29 vdd gnd cell_6t
Xbit_r30_c234 bl_234 br_234 wl_30 vdd gnd cell_6t
Xbit_r31_c234 bl_234 br_234 wl_31 vdd gnd cell_6t
Xbit_r32_c234 bl_234 br_234 wl_32 vdd gnd cell_6t
Xbit_r33_c234 bl_234 br_234 wl_33 vdd gnd cell_6t
Xbit_r34_c234 bl_234 br_234 wl_34 vdd gnd cell_6t
Xbit_r35_c234 bl_234 br_234 wl_35 vdd gnd cell_6t
Xbit_r36_c234 bl_234 br_234 wl_36 vdd gnd cell_6t
Xbit_r37_c234 bl_234 br_234 wl_37 vdd gnd cell_6t
Xbit_r38_c234 bl_234 br_234 wl_38 vdd gnd cell_6t
Xbit_r39_c234 bl_234 br_234 wl_39 vdd gnd cell_6t
Xbit_r40_c234 bl_234 br_234 wl_40 vdd gnd cell_6t
Xbit_r41_c234 bl_234 br_234 wl_41 vdd gnd cell_6t
Xbit_r42_c234 bl_234 br_234 wl_42 vdd gnd cell_6t
Xbit_r43_c234 bl_234 br_234 wl_43 vdd gnd cell_6t
Xbit_r44_c234 bl_234 br_234 wl_44 vdd gnd cell_6t
Xbit_r45_c234 bl_234 br_234 wl_45 vdd gnd cell_6t
Xbit_r46_c234 bl_234 br_234 wl_46 vdd gnd cell_6t
Xbit_r47_c234 bl_234 br_234 wl_47 vdd gnd cell_6t
Xbit_r48_c234 bl_234 br_234 wl_48 vdd gnd cell_6t
Xbit_r49_c234 bl_234 br_234 wl_49 vdd gnd cell_6t
Xbit_r50_c234 bl_234 br_234 wl_50 vdd gnd cell_6t
Xbit_r51_c234 bl_234 br_234 wl_51 vdd gnd cell_6t
Xbit_r52_c234 bl_234 br_234 wl_52 vdd gnd cell_6t
Xbit_r53_c234 bl_234 br_234 wl_53 vdd gnd cell_6t
Xbit_r54_c234 bl_234 br_234 wl_54 vdd gnd cell_6t
Xbit_r55_c234 bl_234 br_234 wl_55 vdd gnd cell_6t
Xbit_r56_c234 bl_234 br_234 wl_56 vdd gnd cell_6t
Xbit_r57_c234 bl_234 br_234 wl_57 vdd gnd cell_6t
Xbit_r58_c234 bl_234 br_234 wl_58 vdd gnd cell_6t
Xbit_r59_c234 bl_234 br_234 wl_59 vdd gnd cell_6t
Xbit_r60_c234 bl_234 br_234 wl_60 vdd gnd cell_6t
Xbit_r61_c234 bl_234 br_234 wl_61 vdd gnd cell_6t
Xbit_r62_c234 bl_234 br_234 wl_62 vdd gnd cell_6t
Xbit_r63_c234 bl_234 br_234 wl_63 vdd gnd cell_6t
Xbit_r64_c234 bl_234 br_234 wl_64 vdd gnd cell_6t
Xbit_r65_c234 bl_234 br_234 wl_65 vdd gnd cell_6t
Xbit_r66_c234 bl_234 br_234 wl_66 vdd gnd cell_6t
Xbit_r67_c234 bl_234 br_234 wl_67 vdd gnd cell_6t
Xbit_r68_c234 bl_234 br_234 wl_68 vdd gnd cell_6t
Xbit_r69_c234 bl_234 br_234 wl_69 vdd gnd cell_6t
Xbit_r70_c234 bl_234 br_234 wl_70 vdd gnd cell_6t
Xbit_r71_c234 bl_234 br_234 wl_71 vdd gnd cell_6t
Xbit_r72_c234 bl_234 br_234 wl_72 vdd gnd cell_6t
Xbit_r73_c234 bl_234 br_234 wl_73 vdd gnd cell_6t
Xbit_r74_c234 bl_234 br_234 wl_74 vdd gnd cell_6t
Xbit_r75_c234 bl_234 br_234 wl_75 vdd gnd cell_6t
Xbit_r76_c234 bl_234 br_234 wl_76 vdd gnd cell_6t
Xbit_r77_c234 bl_234 br_234 wl_77 vdd gnd cell_6t
Xbit_r78_c234 bl_234 br_234 wl_78 vdd gnd cell_6t
Xbit_r79_c234 bl_234 br_234 wl_79 vdd gnd cell_6t
Xbit_r80_c234 bl_234 br_234 wl_80 vdd gnd cell_6t
Xbit_r81_c234 bl_234 br_234 wl_81 vdd gnd cell_6t
Xbit_r82_c234 bl_234 br_234 wl_82 vdd gnd cell_6t
Xbit_r83_c234 bl_234 br_234 wl_83 vdd gnd cell_6t
Xbit_r84_c234 bl_234 br_234 wl_84 vdd gnd cell_6t
Xbit_r85_c234 bl_234 br_234 wl_85 vdd gnd cell_6t
Xbit_r86_c234 bl_234 br_234 wl_86 vdd gnd cell_6t
Xbit_r87_c234 bl_234 br_234 wl_87 vdd gnd cell_6t
Xbit_r88_c234 bl_234 br_234 wl_88 vdd gnd cell_6t
Xbit_r89_c234 bl_234 br_234 wl_89 vdd gnd cell_6t
Xbit_r90_c234 bl_234 br_234 wl_90 vdd gnd cell_6t
Xbit_r91_c234 bl_234 br_234 wl_91 vdd gnd cell_6t
Xbit_r92_c234 bl_234 br_234 wl_92 vdd gnd cell_6t
Xbit_r93_c234 bl_234 br_234 wl_93 vdd gnd cell_6t
Xbit_r94_c234 bl_234 br_234 wl_94 vdd gnd cell_6t
Xbit_r95_c234 bl_234 br_234 wl_95 vdd gnd cell_6t
Xbit_r96_c234 bl_234 br_234 wl_96 vdd gnd cell_6t
Xbit_r97_c234 bl_234 br_234 wl_97 vdd gnd cell_6t
Xbit_r98_c234 bl_234 br_234 wl_98 vdd gnd cell_6t
Xbit_r99_c234 bl_234 br_234 wl_99 vdd gnd cell_6t
Xbit_r100_c234 bl_234 br_234 wl_100 vdd gnd cell_6t
Xbit_r101_c234 bl_234 br_234 wl_101 vdd gnd cell_6t
Xbit_r102_c234 bl_234 br_234 wl_102 vdd gnd cell_6t
Xbit_r103_c234 bl_234 br_234 wl_103 vdd gnd cell_6t
Xbit_r104_c234 bl_234 br_234 wl_104 vdd gnd cell_6t
Xbit_r105_c234 bl_234 br_234 wl_105 vdd gnd cell_6t
Xbit_r106_c234 bl_234 br_234 wl_106 vdd gnd cell_6t
Xbit_r107_c234 bl_234 br_234 wl_107 vdd gnd cell_6t
Xbit_r108_c234 bl_234 br_234 wl_108 vdd gnd cell_6t
Xbit_r109_c234 bl_234 br_234 wl_109 vdd gnd cell_6t
Xbit_r110_c234 bl_234 br_234 wl_110 vdd gnd cell_6t
Xbit_r111_c234 bl_234 br_234 wl_111 vdd gnd cell_6t
Xbit_r112_c234 bl_234 br_234 wl_112 vdd gnd cell_6t
Xbit_r113_c234 bl_234 br_234 wl_113 vdd gnd cell_6t
Xbit_r114_c234 bl_234 br_234 wl_114 vdd gnd cell_6t
Xbit_r115_c234 bl_234 br_234 wl_115 vdd gnd cell_6t
Xbit_r116_c234 bl_234 br_234 wl_116 vdd gnd cell_6t
Xbit_r117_c234 bl_234 br_234 wl_117 vdd gnd cell_6t
Xbit_r118_c234 bl_234 br_234 wl_118 vdd gnd cell_6t
Xbit_r119_c234 bl_234 br_234 wl_119 vdd gnd cell_6t
Xbit_r120_c234 bl_234 br_234 wl_120 vdd gnd cell_6t
Xbit_r121_c234 bl_234 br_234 wl_121 vdd gnd cell_6t
Xbit_r122_c234 bl_234 br_234 wl_122 vdd gnd cell_6t
Xbit_r123_c234 bl_234 br_234 wl_123 vdd gnd cell_6t
Xbit_r124_c234 bl_234 br_234 wl_124 vdd gnd cell_6t
Xbit_r125_c234 bl_234 br_234 wl_125 vdd gnd cell_6t
Xbit_r126_c234 bl_234 br_234 wl_126 vdd gnd cell_6t
Xbit_r127_c234 bl_234 br_234 wl_127 vdd gnd cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd cell_6t
Xbit_r1_c235 bl_235 br_235 wl_1 vdd gnd cell_6t
Xbit_r2_c235 bl_235 br_235 wl_2 vdd gnd cell_6t
Xbit_r3_c235 bl_235 br_235 wl_3 vdd gnd cell_6t
Xbit_r4_c235 bl_235 br_235 wl_4 vdd gnd cell_6t
Xbit_r5_c235 bl_235 br_235 wl_5 vdd gnd cell_6t
Xbit_r6_c235 bl_235 br_235 wl_6 vdd gnd cell_6t
Xbit_r7_c235 bl_235 br_235 wl_7 vdd gnd cell_6t
Xbit_r8_c235 bl_235 br_235 wl_8 vdd gnd cell_6t
Xbit_r9_c235 bl_235 br_235 wl_9 vdd gnd cell_6t
Xbit_r10_c235 bl_235 br_235 wl_10 vdd gnd cell_6t
Xbit_r11_c235 bl_235 br_235 wl_11 vdd gnd cell_6t
Xbit_r12_c235 bl_235 br_235 wl_12 vdd gnd cell_6t
Xbit_r13_c235 bl_235 br_235 wl_13 vdd gnd cell_6t
Xbit_r14_c235 bl_235 br_235 wl_14 vdd gnd cell_6t
Xbit_r15_c235 bl_235 br_235 wl_15 vdd gnd cell_6t
Xbit_r16_c235 bl_235 br_235 wl_16 vdd gnd cell_6t
Xbit_r17_c235 bl_235 br_235 wl_17 vdd gnd cell_6t
Xbit_r18_c235 bl_235 br_235 wl_18 vdd gnd cell_6t
Xbit_r19_c235 bl_235 br_235 wl_19 vdd gnd cell_6t
Xbit_r20_c235 bl_235 br_235 wl_20 vdd gnd cell_6t
Xbit_r21_c235 bl_235 br_235 wl_21 vdd gnd cell_6t
Xbit_r22_c235 bl_235 br_235 wl_22 vdd gnd cell_6t
Xbit_r23_c235 bl_235 br_235 wl_23 vdd gnd cell_6t
Xbit_r24_c235 bl_235 br_235 wl_24 vdd gnd cell_6t
Xbit_r25_c235 bl_235 br_235 wl_25 vdd gnd cell_6t
Xbit_r26_c235 bl_235 br_235 wl_26 vdd gnd cell_6t
Xbit_r27_c235 bl_235 br_235 wl_27 vdd gnd cell_6t
Xbit_r28_c235 bl_235 br_235 wl_28 vdd gnd cell_6t
Xbit_r29_c235 bl_235 br_235 wl_29 vdd gnd cell_6t
Xbit_r30_c235 bl_235 br_235 wl_30 vdd gnd cell_6t
Xbit_r31_c235 bl_235 br_235 wl_31 vdd gnd cell_6t
Xbit_r32_c235 bl_235 br_235 wl_32 vdd gnd cell_6t
Xbit_r33_c235 bl_235 br_235 wl_33 vdd gnd cell_6t
Xbit_r34_c235 bl_235 br_235 wl_34 vdd gnd cell_6t
Xbit_r35_c235 bl_235 br_235 wl_35 vdd gnd cell_6t
Xbit_r36_c235 bl_235 br_235 wl_36 vdd gnd cell_6t
Xbit_r37_c235 bl_235 br_235 wl_37 vdd gnd cell_6t
Xbit_r38_c235 bl_235 br_235 wl_38 vdd gnd cell_6t
Xbit_r39_c235 bl_235 br_235 wl_39 vdd gnd cell_6t
Xbit_r40_c235 bl_235 br_235 wl_40 vdd gnd cell_6t
Xbit_r41_c235 bl_235 br_235 wl_41 vdd gnd cell_6t
Xbit_r42_c235 bl_235 br_235 wl_42 vdd gnd cell_6t
Xbit_r43_c235 bl_235 br_235 wl_43 vdd gnd cell_6t
Xbit_r44_c235 bl_235 br_235 wl_44 vdd gnd cell_6t
Xbit_r45_c235 bl_235 br_235 wl_45 vdd gnd cell_6t
Xbit_r46_c235 bl_235 br_235 wl_46 vdd gnd cell_6t
Xbit_r47_c235 bl_235 br_235 wl_47 vdd gnd cell_6t
Xbit_r48_c235 bl_235 br_235 wl_48 vdd gnd cell_6t
Xbit_r49_c235 bl_235 br_235 wl_49 vdd gnd cell_6t
Xbit_r50_c235 bl_235 br_235 wl_50 vdd gnd cell_6t
Xbit_r51_c235 bl_235 br_235 wl_51 vdd gnd cell_6t
Xbit_r52_c235 bl_235 br_235 wl_52 vdd gnd cell_6t
Xbit_r53_c235 bl_235 br_235 wl_53 vdd gnd cell_6t
Xbit_r54_c235 bl_235 br_235 wl_54 vdd gnd cell_6t
Xbit_r55_c235 bl_235 br_235 wl_55 vdd gnd cell_6t
Xbit_r56_c235 bl_235 br_235 wl_56 vdd gnd cell_6t
Xbit_r57_c235 bl_235 br_235 wl_57 vdd gnd cell_6t
Xbit_r58_c235 bl_235 br_235 wl_58 vdd gnd cell_6t
Xbit_r59_c235 bl_235 br_235 wl_59 vdd gnd cell_6t
Xbit_r60_c235 bl_235 br_235 wl_60 vdd gnd cell_6t
Xbit_r61_c235 bl_235 br_235 wl_61 vdd gnd cell_6t
Xbit_r62_c235 bl_235 br_235 wl_62 vdd gnd cell_6t
Xbit_r63_c235 bl_235 br_235 wl_63 vdd gnd cell_6t
Xbit_r64_c235 bl_235 br_235 wl_64 vdd gnd cell_6t
Xbit_r65_c235 bl_235 br_235 wl_65 vdd gnd cell_6t
Xbit_r66_c235 bl_235 br_235 wl_66 vdd gnd cell_6t
Xbit_r67_c235 bl_235 br_235 wl_67 vdd gnd cell_6t
Xbit_r68_c235 bl_235 br_235 wl_68 vdd gnd cell_6t
Xbit_r69_c235 bl_235 br_235 wl_69 vdd gnd cell_6t
Xbit_r70_c235 bl_235 br_235 wl_70 vdd gnd cell_6t
Xbit_r71_c235 bl_235 br_235 wl_71 vdd gnd cell_6t
Xbit_r72_c235 bl_235 br_235 wl_72 vdd gnd cell_6t
Xbit_r73_c235 bl_235 br_235 wl_73 vdd gnd cell_6t
Xbit_r74_c235 bl_235 br_235 wl_74 vdd gnd cell_6t
Xbit_r75_c235 bl_235 br_235 wl_75 vdd gnd cell_6t
Xbit_r76_c235 bl_235 br_235 wl_76 vdd gnd cell_6t
Xbit_r77_c235 bl_235 br_235 wl_77 vdd gnd cell_6t
Xbit_r78_c235 bl_235 br_235 wl_78 vdd gnd cell_6t
Xbit_r79_c235 bl_235 br_235 wl_79 vdd gnd cell_6t
Xbit_r80_c235 bl_235 br_235 wl_80 vdd gnd cell_6t
Xbit_r81_c235 bl_235 br_235 wl_81 vdd gnd cell_6t
Xbit_r82_c235 bl_235 br_235 wl_82 vdd gnd cell_6t
Xbit_r83_c235 bl_235 br_235 wl_83 vdd gnd cell_6t
Xbit_r84_c235 bl_235 br_235 wl_84 vdd gnd cell_6t
Xbit_r85_c235 bl_235 br_235 wl_85 vdd gnd cell_6t
Xbit_r86_c235 bl_235 br_235 wl_86 vdd gnd cell_6t
Xbit_r87_c235 bl_235 br_235 wl_87 vdd gnd cell_6t
Xbit_r88_c235 bl_235 br_235 wl_88 vdd gnd cell_6t
Xbit_r89_c235 bl_235 br_235 wl_89 vdd gnd cell_6t
Xbit_r90_c235 bl_235 br_235 wl_90 vdd gnd cell_6t
Xbit_r91_c235 bl_235 br_235 wl_91 vdd gnd cell_6t
Xbit_r92_c235 bl_235 br_235 wl_92 vdd gnd cell_6t
Xbit_r93_c235 bl_235 br_235 wl_93 vdd gnd cell_6t
Xbit_r94_c235 bl_235 br_235 wl_94 vdd gnd cell_6t
Xbit_r95_c235 bl_235 br_235 wl_95 vdd gnd cell_6t
Xbit_r96_c235 bl_235 br_235 wl_96 vdd gnd cell_6t
Xbit_r97_c235 bl_235 br_235 wl_97 vdd gnd cell_6t
Xbit_r98_c235 bl_235 br_235 wl_98 vdd gnd cell_6t
Xbit_r99_c235 bl_235 br_235 wl_99 vdd gnd cell_6t
Xbit_r100_c235 bl_235 br_235 wl_100 vdd gnd cell_6t
Xbit_r101_c235 bl_235 br_235 wl_101 vdd gnd cell_6t
Xbit_r102_c235 bl_235 br_235 wl_102 vdd gnd cell_6t
Xbit_r103_c235 bl_235 br_235 wl_103 vdd gnd cell_6t
Xbit_r104_c235 bl_235 br_235 wl_104 vdd gnd cell_6t
Xbit_r105_c235 bl_235 br_235 wl_105 vdd gnd cell_6t
Xbit_r106_c235 bl_235 br_235 wl_106 vdd gnd cell_6t
Xbit_r107_c235 bl_235 br_235 wl_107 vdd gnd cell_6t
Xbit_r108_c235 bl_235 br_235 wl_108 vdd gnd cell_6t
Xbit_r109_c235 bl_235 br_235 wl_109 vdd gnd cell_6t
Xbit_r110_c235 bl_235 br_235 wl_110 vdd gnd cell_6t
Xbit_r111_c235 bl_235 br_235 wl_111 vdd gnd cell_6t
Xbit_r112_c235 bl_235 br_235 wl_112 vdd gnd cell_6t
Xbit_r113_c235 bl_235 br_235 wl_113 vdd gnd cell_6t
Xbit_r114_c235 bl_235 br_235 wl_114 vdd gnd cell_6t
Xbit_r115_c235 bl_235 br_235 wl_115 vdd gnd cell_6t
Xbit_r116_c235 bl_235 br_235 wl_116 vdd gnd cell_6t
Xbit_r117_c235 bl_235 br_235 wl_117 vdd gnd cell_6t
Xbit_r118_c235 bl_235 br_235 wl_118 vdd gnd cell_6t
Xbit_r119_c235 bl_235 br_235 wl_119 vdd gnd cell_6t
Xbit_r120_c235 bl_235 br_235 wl_120 vdd gnd cell_6t
Xbit_r121_c235 bl_235 br_235 wl_121 vdd gnd cell_6t
Xbit_r122_c235 bl_235 br_235 wl_122 vdd gnd cell_6t
Xbit_r123_c235 bl_235 br_235 wl_123 vdd gnd cell_6t
Xbit_r124_c235 bl_235 br_235 wl_124 vdd gnd cell_6t
Xbit_r125_c235 bl_235 br_235 wl_125 vdd gnd cell_6t
Xbit_r126_c235 bl_235 br_235 wl_126 vdd gnd cell_6t
Xbit_r127_c235 bl_235 br_235 wl_127 vdd gnd cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd cell_6t
Xbit_r1_c236 bl_236 br_236 wl_1 vdd gnd cell_6t
Xbit_r2_c236 bl_236 br_236 wl_2 vdd gnd cell_6t
Xbit_r3_c236 bl_236 br_236 wl_3 vdd gnd cell_6t
Xbit_r4_c236 bl_236 br_236 wl_4 vdd gnd cell_6t
Xbit_r5_c236 bl_236 br_236 wl_5 vdd gnd cell_6t
Xbit_r6_c236 bl_236 br_236 wl_6 vdd gnd cell_6t
Xbit_r7_c236 bl_236 br_236 wl_7 vdd gnd cell_6t
Xbit_r8_c236 bl_236 br_236 wl_8 vdd gnd cell_6t
Xbit_r9_c236 bl_236 br_236 wl_9 vdd gnd cell_6t
Xbit_r10_c236 bl_236 br_236 wl_10 vdd gnd cell_6t
Xbit_r11_c236 bl_236 br_236 wl_11 vdd gnd cell_6t
Xbit_r12_c236 bl_236 br_236 wl_12 vdd gnd cell_6t
Xbit_r13_c236 bl_236 br_236 wl_13 vdd gnd cell_6t
Xbit_r14_c236 bl_236 br_236 wl_14 vdd gnd cell_6t
Xbit_r15_c236 bl_236 br_236 wl_15 vdd gnd cell_6t
Xbit_r16_c236 bl_236 br_236 wl_16 vdd gnd cell_6t
Xbit_r17_c236 bl_236 br_236 wl_17 vdd gnd cell_6t
Xbit_r18_c236 bl_236 br_236 wl_18 vdd gnd cell_6t
Xbit_r19_c236 bl_236 br_236 wl_19 vdd gnd cell_6t
Xbit_r20_c236 bl_236 br_236 wl_20 vdd gnd cell_6t
Xbit_r21_c236 bl_236 br_236 wl_21 vdd gnd cell_6t
Xbit_r22_c236 bl_236 br_236 wl_22 vdd gnd cell_6t
Xbit_r23_c236 bl_236 br_236 wl_23 vdd gnd cell_6t
Xbit_r24_c236 bl_236 br_236 wl_24 vdd gnd cell_6t
Xbit_r25_c236 bl_236 br_236 wl_25 vdd gnd cell_6t
Xbit_r26_c236 bl_236 br_236 wl_26 vdd gnd cell_6t
Xbit_r27_c236 bl_236 br_236 wl_27 vdd gnd cell_6t
Xbit_r28_c236 bl_236 br_236 wl_28 vdd gnd cell_6t
Xbit_r29_c236 bl_236 br_236 wl_29 vdd gnd cell_6t
Xbit_r30_c236 bl_236 br_236 wl_30 vdd gnd cell_6t
Xbit_r31_c236 bl_236 br_236 wl_31 vdd gnd cell_6t
Xbit_r32_c236 bl_236 br_236 wl_32 vdd gnd cell_6t
Xbit_r33_c236 bl_236 br_236 wl_33 vdd gnd cell_6t
Xbit_r34_c236 bl_236 br_236 wl_34 vdd gnd cell_6t
Xbit_r35_c236 bl_236 br_236 wl_35 vdd gnd cell_6t
Xbit_r36_c236 bl_236 br_236 wl_36 vdd gnd cell_6t
Xbit_r37_c236 bl_236 br_236 wl_37 vdd gnd cell_6t
Xbit_r38_c236 bl_236 br_236 wl_38 vdd gnd cell_6t
Xbit_r39_c236 bl_236 br_236 wl_39 vdd gnd cell_6t
Xbit_r40_c236 bl_236 br_236 wl_40 vdd gnd cell_6t
Xbit_r41_c236 bl_236 br_236 wl_41 vdd gnd cell_6t
Xbit_r42_c236 bl_236 br_236 wl_42 vdd gnd cell_6t
Xbit_r43_c236 bl_236 br_236 wl_43 vdd gnd cell_6t
Xbit_r44_c236 bl_236 br_236 wl_44 vdd gnd cell_6t
Xbit_r45_c236 bl_236 br_236 wl_45 vdd gnd cell_6t
Xbit_r46_c236 bl_236 br_236 wl_46 vdd gnd cell_6t
Xbit_r47_c236 bl_236 br_236 wl_47 vdd gnd cell_6t
Xbit_r48_c236 bl_236 br_236 wl_48 vdd gnd cell_6t
Xbit_r49_c236 bl_236 br_236 wl_49 vdd gnd cell_6t
Xbit_r50_c236 bl_236 br_236 wl_50 vdd gnd cell_6t
Xbit_r51_c236 bl_236 br_236 wl_51 vdd gnd cell_6t
Xbit_r52_c236 bl_236 br_236 wl_52 vdd gnd cell_6t
Xbit_r53_c236 bl_236 br_236 wl_53 vdd gnd cell_6t
Xbit_r54_c236 bl_236 br_236 wl_54 vdd gnd cell_6t
Xbit_r55_c236 bl_236 br_236 wl_55 vdd gnd cell_6t
Xbit_r56_c236 bl_236 br_236 wl_56 vdd gnd cell_6t
Xbit_r57_c236 bl_236 br_236 wl_57 vdd gnd cell_6t
Xbit_r58_c236 bl_236 br_236 wl_58 vdd gnd cell_6t
Xbit_r59_c236 bl_236 br_236 wl_59 vdd gnd cell_6t
Xbit_r60_c236 bl_236 br_236 wl_60 vdd gnd cell_6t
Xbit_r61_c236 bl_236 br_236 wl_61 vdd gnd cell_6t
Xbit_r62_c236 bl_236 br_236 wl_62 vdd gnd cell_6t
Xbit_r63_c236 bl_236 br_236 wl_63 vdd gnd cell_6t
Xbit_r64_c236 bl_236 br_236 wl_64 vdd gnd cell_6t
Xbit_r65_c236 bl_236 br_236 wl_65 vdd gnd cell_6t
Xbit_r66_c236 bl_236 br_236 wl_66 vdd gnd cell_6t
Xbit_r67_c236 bl_236 br_236 wl_67 vdd gnd cell_6t
Xbit_r68_c236 bl_236 br_236 wl_68 vdd gnd cell_6t
Xbit_r69_c236 bl_236 br_236 wl_69 vdd gnd cell_6t
Xbit_r70_c236 bl_236 br_236 wl_70 vdd gnd cell_6t
Xbit_r71_c236 bl_236 br_236 wl_71 vdd gnd cell_6t
Xbit_r72_c236 bl_236 br_236 wl_72 vdd gnd cell_6t
Xbit_r73_c236 bl_236 br_236 wl_73 vdd gnd cell_6t
Xbit_r74_c236 bl_236 br_236 wl_74 vdd gnd cell_6t
Xbit_r75_c236 bl_236 br_236 wl_75 vdd gnd cell_6t
Xbit_r76_c236 bl_236 br_236 wl_76 vdd gnd cell_6t
Xbit_r77_c236 bl_236 br_236 wl_77 vdd gnd cell_6t
Xbit_r78_c236 bl_236 br_236 wl_78 vdd gnd cell_6t
Xbit_r79_c236 bl_236 br_236 wl_79 vdd gnd cell_6t
Xbit_r80_c236 bl_236 br_236 wl_80 vdd gnd cell_6t
Xbit_r81_c236 bl_236 br_236 wl_81 vdd gnd cell_6t
Xbit_r82_c236 bl_236 br_236 wl_82 vdd gnd cell_6t
Xbit_r83_c236 bl_236 br_236 wl_83 vdd gnd cell_6t
Xbit_r84_c236 bl_236 br_236 wl_84 vdd gnd cell_6t
Xbit_r85_c236 bl_236 br_236 wl_85 vdd gnd cell_6t
Xbit_r86_c236 bl_236 br_236 wl_86 vdd gnd cell_6t
Xbit_r87_c236 bl_236 br_236 wl_87 vdd gnd cell_6t
Xbit_r88_c236 bl_236 br_236 wl_88 vdd gnd cell_6t
Xbit_r89_c236 bl_236 br_236 wl_89 vdd gnd cell_6t
Xbit_r90_c236 bl_236 br_236 wl_90 vdd gnd cell_6t
Xbit_r91_c236 bl_236 br_236 wl_91 vdd gnd cell_6t
Xbit_r92_c236 bl_236 br_236 wl_92 vdd gnd cell_6t
Xbit_r93_c236 bl_236 br_236 wl_93 vdd gnd cell_6t
Xbit_r94_c236 bl_236 br_236 wl_94 vdd gnd cell_6t
Xbit_r95_c236 bl_236 br_236 wl_95 vdd gnd cell_6t
Xbit_r96_c236 bl_236 br_236 wl_96 vdd gnd cell_6t
Xbit_r97_c236 bl_236 br_236 wl_97 vdd gnd cell_6t
Xbit_r98_c236 bl_236 br_236 wl_98 vdd gnd cell_6t
Xbit_r99_c236 bl_236 br_236 wl_99 vdd gnd cell_6t
Xbit_r100_c236 bl_236 br_236 wl_100 vdd gnd cell_6t
Xbit_r101_c236 bl_236 br_236 wl_101 vdd gnd cell_6t
Xbit_r102_c236 bl_236 br_236 wl_102 vdd gnd cell_6t
Xbit_r103_c236 bl_236 br_236 wl_103 vdd gnd cell_6t
Xbit_r104_c236 bl_236 br_236 wl_104 vdd gnd cell_6t
Xbit_r105_c236 bl_236 br_236 wl_105 vdd gnd cell_6t
Xbit_r106_c236 bl_236 br_236 wl_106 vdd gnd cell_6t
Xbit_r107_c236 bl_236 br_236 wl_107 vdd gnd cell_6t
Xbit_r108_c236 bl_236 br_236 wl_108 vdd gnd cell_6t
Xbit_r109_c236 bl_236 br_236 wl_109 vdd gnd cell_6t
Xbit_r110_c236 bl_236 br_236 wl_110 vdd gnd cell_6t
Xbit_r111_c236 bl_236 br_236 wl_111 vdd gnd cell_6t
Xbit_r112_c236 bl_236 br_236 wl_112 vdd gnd cell_6t
Xbit_r113_c236 bl_236 br_236 wl_113 vdd gnd cell_6t
Xbit_r114_c236 bl_236 br_236 wl_114 vdd gnd cell_6t
Xbit_r115_c236 bl_236 br_236 wl_115 vdd gnd cell_6t
Xbit_r116_c236 bl_236 br_236 wl_116 vdd gnd cell_6t
Xbit_r117_c236 bl_236 br_236 wl_117 vdd gnd cell_6t
Xbit_r118_c236 bl_236 br_236 wl_118 vdd gnd cell_6t
Xbit_r119_c236 bl_236 br_236 wl_119 vdd gnd cell_6t
Xbit_r120_c236 bl_236 br_236 wl_120 vdd gnd cell_6t
Xbit_r121_c236 bl_236 br_236 wl_121 vdd gnd cell_6t
Xbit_r122_c236 bl_236 br_236 wl_122 vdd gnd cell_6t
Xbit_r123_c236 bl_236 br_236 wl_123 vdd gnd cell_6t
Xbit_r124_c236 bl_236 br_236 wl_124 vdd gnd cell_6t
Xbit_r125_c236 bl_236 br_236 wl_125 vdd gnd cell_6t
Xbit_r126_c236 bl_236 br_236 wl_126 vdd gnd cell_6t
Xbit_r127_c236 bl_236 br_236 wl_127 vdd gnd cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd cell_6t
Xbit_r1_c237 bl_237 br_237 wl_1 vdd gnd cell_6t
Xbit_r2_c237 bl_237 br_237 wl_2 vdd gnd cell_6t
Xbit_r3_c237 bl_237 br_237 wl_3 vdd gnd cell_6t
Xbit_r4_c237 bl_237 br_237 wl_4 vdd gnd cell_6t
Xbit_r5_c237 bl_237 br_237 wl_5 vdd gnd cell_6t
Xbit_r6_c237 bl_237 br_237 wl_6 vdd gnd cell_6t
Xbit_r7_c237 bl_237 br_237 wl_7 vdd gnd cell_6t
Xbit_r8_c237 bl_237 br_237 wl_8 vdd gnd cell_6t
Xbit_r9_c237 bl_237 br_237 wl_9 vdd gnd cell_6t
Xbit_r10_c237 bl_237 br_237 wl_10 vdd gnd cell_6t
Xbit_r11_c237 bl_237 br_237 wl_11 vdd gnd cell_6t
Xbit_r12_c237 bl_237 br_237 wl_12 vdd gnd cell_6t
Xbit_r13_c237 bl_237 br_237 wl_13 vdd gnd cell_6t
Xbit_r14_c237 bl_237 br_237 wl_14 vdd gnd cell_6t
Xbit_r15_c237 bl_237 br_237 wl_15 vdd gnd cell_6t
Xbit_r16_c237 bl_237 br_237 wl_16 vdd gnd cell_6t
Xbit_r17_c237 bl_237 br_237 wl_17 vdd gnd cell_6t
Xbit_r18_c237 bl_237 br_237 wl_18 vdd gnd cell_6t
Xbit_r19_c237 bl_237 br_237 wl_19 vdd gnd cell_6t
Xbit_r20_c237 bl_237 br_237 wl_20 vdd gnd cell_6t
Xbit_r21_c237 bl_237 br_237 wl_21 vdd gnd cell_6t
Xbit_r22_c237 bl_237 br_237 wl_22 vdd gnd cell_6t
Xbit_r23_c237 bl_237 br_237 wl_23 vdd gnd cell_6t
Xbit_r24_c237 bl_237 br_237 wl_24 vdd gnd cell_6t
Xbit_r25_c237 bl_237 br_237 wl_25 vdd gnd cell_6t
Xbit_r26_c237 bl_237 br_237 wl_26 vdd gnd cell_6t
Xbit_r27_c237 bl_237 br_237 wl_27 vdd gnd cell_6t
Xbit_r28_c237 bl_237 br_237 wl_28 vdd gnd cell_6t
Xbit_r29_c237 bl_237 br_237 wl_29 vdd gnd cell_6t
Xbit_r30_c237 bl_237 br_237 wl_30 vdd gnd cell_6t
Xbit_r31_c237 bl_237 br_237 wl_31 vdd gnd cell_6t
Xbit_r32_c237 bl_237 br_237 wl_32 vdd gnd cell_6t
Xbit_r33_c237 bl_237 br_237 wl_33 vdd gnd cell_6t
Xbit_r34_c237 bl_237 br_237 wl_34 vdd gnd cell_6t
Xbit_r35_c237 bl_237 br_237 wl_35 vdd gnd cell_6t
Xbit_r36_c237 bl_237 br_237 wl_36 vdd gnd cell_6t
Xbit_r37_c237 bl_237 br_237 wl_37 vdd gnd cell_6t
Xbit_r38_c237 bl_237 br_237 wl_38 vdd gnd cell_6t
Xbit_r39_c237 bl_237 br_237 wl_39 vdd gnd cell_6t
Xbit_r40_c237 bl_237 br_237 wl_40 vdd gnd cell_6t
Xbit_r41_c237 bl_237 br_237 wl_41 vdd gnd cell_6t
Xbit_r42_c237 bl_237 br_237 wl_42 vdd gnd cell_6t
Xbit_r43_c237 bl_237 br_237 wl_43 vdd gnd cell_6t
Xbit_r44_c237 bl_237 br_237 wl_44 vdd gnd cell_6t
Xbit_r45_c237 bl_237 br_237 wl_45 vdd gnd cell_6t
Xbit_r46_c237 bl_237 br_237 wl_46 vdd gnd cell_6t
Xbit_r47_c237 bl_237 br_237 wl_47 vdd gnd cell_6t
Xbit_r48_c237 bl_237 br_237 wl_48 vdd gnd cell_6t
Xbit_r49_c237 bl_237 br_237 wl_49 vdd gnd cell_6t
Xbit_r50_c237 bl_237 br_237 wl_50 vdd gnd cell_6t
Xbit_r51_c237 bl_237 br_237 wl_51 vdd gnd cell_6t
Xbit_r52_c237 bl_237 br_237 wl_52 vdd gnd cell_6t
Xbit_r53_c237 bl_237 br_237 wl_53 vdd gnd cell_6t
Xbit_r54_c237 bl_237 br_237 wl_54 vdd gnd cell_6t
Xbit_r55_c237 bl_237 br_237 wl_55 vdd gnd cell_6t
Xbit_r56_c237 bl_237 br_237 wl_56 vdd gnd cell_6t
Xbit_r57_c237 bl_237 br_237 wl_57 vdd gnd cell_6t
Xbit_r58_c237 bl_237 br_237 wl_58 vdd gnd cell_6t
Xbit_r59_c237 bl_237 br_237 wl_59 vdd gnd cell_6t
Xbit_r60_c237 bl_237 br_237 wl_60 vdd gnd cell_6t
Xbit_r61_c237 bl_237 br_237 wl_61 vdd gnd cell_6t
Xbit_r62_c237 bl_237 br_237 wl_62 vdd gnd cell_6t
Xbit_r63_c237 bl_237 br_237 wl_63 vdd gnd cell_6t
Xbit_r64_c237 bl_237 br_237 wl_64 vdd gnd cell_6t
Xbit_r65_c237 bl_237 br_237 wl_65 vdd gnd cell_6t
Xbit_r66_c237 bl_237 br_237 wl_66 vdd gnd cell_6t
Xbit_r67_c237 bl_237 br_237 wl_67 vdd gnd cell_6t
Xbit_r68_c237 bl_237 br_237 wl_68 vdd gnd cell_6t
Xbit_r69_c237 bl_237 br_237 wl_69 vdd gnd cell_6t
Xbit_r70_c237 bl_237 br_237 wl_70 vdd gnd cell_6t
Xbit_r71_c237 bl_237 br_237 wl_71 vdd gnd cell_6t
Xbit_r72_c237 bl_237 br_237 wl_72 vdd gnd cell_6t
Xbit_r73_c237 bl_237 br_237 wl_73 vdd gnd cell_6t
Xbit_r74_c237 bl_237 br_237 wl_74 vdd gnd cell_6t
Xbit_r75_c237 bl_237 br_237 wl_75 vdd gnd cell_6t
Xbit_r76_c237 bl_237 br_237 wl_76 vdd gnd cell_6t
Xbit_r77_c237 bl_237 br_237 wl_77 vdd gnd cell_6t
Xbit_r78_c237 bl_237 br_237 wl_78 vdd gnd cell_6t
Xbit_r79_c237 bl_237 br_237 wl_79 vdd gnd cell_6t
Xbit_r80_c237 bl_237 br_237 wl_80 vdd gnd cell_6t
Xbit_r81_c237 bl_237 br_237 wl_81 vdd gnd cell_6t
Xbit_r82_c237 bl_237 br_237 wl_82 vdd gnd cell_6t
Xbit_r83_c237 bl_237 br_237 wl_83 vdd gnd cell_6t
Xbit_r84_c237 bl_237 br_237 wl_84 vdd gnd cell_6t
Xbit_r85_c237 bl_237 br_237 wl_85 vdd gnd cell_6t
Xbit_r86_c237 bl_237 br_237 wl_86 vdd gnd cell_6t
Xbit_r87_c237 bl_237 br_237 wl_87 vdd gnd cell_6t
Xbit_r88_c237 bl_237 br_237 wl_88 vdd gnd cell_6t
Xbit_r89_c237 bl_237 br_237 wl_89 vdd gnd cell_6t
Xbit_r90_c237 bl_237 br_237 wl_90 vdd gnd cell_6t
Xbit_r91_c237 bl_237 br_237 wl_91 vdd gnd cell_6t
Xbit_r92_c237 bl_237 br_237 wl_92 vdd gnd cell_6t
Xbit_r93_c237 bl_237 br_237 wl_93 vdd gnd cell_6t
Xbit_r94_c237 bl_237 br_237 wl_94 vdd gnd cell_6t
Xbit_r95_c237 bl_237 br_237 wl_95 vdd gnd cell_6t
Xbit_r96_c237 bl_237 br_237 wl_96 vdd gnd cell_6t
Xbit_r97_c237 bl_237 br_237 wl_97 vdd gnd cell_6t
Xbit_r98_c237 bl_237 br_237 wl_98 vdd gnd cell_6t
Xbit_r99_c237 bl_237 br_237 wl_99 vdd gnd cell_6t
Xbit_r100_c237 bl_237 br_237 wl_100 vdd gnd cell_6t
Xbit_r101_c237 bl_237 br_237 wl_101 vdd gnd cell_6t
Xbit_r102_c237 bl_237 br_237 wl_102 vdd gnd cell_6t
Xbit_r103_c237 bl_237 br_237 wl_103 vdd gnd cell_6t
Xbit_r104_c237 bl_237 br_237 wl_104 vdd gnd cell_6t
Xbit_r105_c237 bl_237 br_237 wl_105 vdd gnd cell_6t
Xbit_r106_c237 bl_237 br_237 wl_106 vdd gnd cell_6t
Xbit_r107_c237 bl_237 br_237 wl_107 vdd gnd cell_6t
Xbit_r108_c237 bl_237 br_237 wl_108 vdd gnd cell_6t
Xbit_r109_c237 bl_237 br_237 wl_109 vdd gnd cell_6t
Xbit_r110_c237 bl_237 br_237 wl_110 vdd gnd cell_6t
Xbit_r111_c237 bl_237 br_237 wl_111 vdd gnd cell_6t
Xbit_r112_c237 bl_237 br_237 wl_112 vdd gnd cell_6t
Xbit_r113_c237 bl_237 br_237 wl_113 vdd gnd cell_6t
Xbit_r114_c237 bl_237 br_237 wl_114 vdd gnd cell_6t
Xbit_r115_c237 bl_237 br_237 wl_115 vdd gnd cell_6t
Xbit_r116_c237 bl_237 br_237 wl_116 vdd gnd cell_6t
Xbit_r117_c237 bl_237 br_237 wl_117 vdd gnd cell_6t
Xbit_r118_c237 bl_237 br_237 wl_118 vdd gnd cell_6t
Xbit_r119_c237 bl_237 br_237 wl_119 vdd gnd cell_6t
Xbit_r120_c237 bl_237 br_237 wl_120 vdd gnd cell_6t
Xbit_r121_c237 bl_237 br_237 wl_121 vdd gnd cell_6t
Xbit_r122_c237 bl_237 br_237 wl_122 vdd gnd cell_6t
Xbit_r123_c237 bl_237 br_237 wl_123 vdd gnd cell_6t
Xbit_r124_c237 bl_237 br_237 wl_124 vdd gnd cell_6t
Xbit_r125_c237 bl_237 br_237 wl_125 vdd gnd cell_6t
Xbit_r126_c237 bl_237 br_237 wl_126 vdd gnd cell_6t
Xbit_r127_c237 bl_237 br_237 wl_127 vdd gnd cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd cell_6t
Xbit_r1_c238 bl_238 br_238 wl_1 vdd gnd cell_6t
Xbit_r2_c238 bl_238 br_238 wl_2 vdd gnd cell_6t
Xbit_r3_c238 bl_238 br_238 wl_3 vdd gnd cell_6t
Xbit_r4_c238 bl_238 br_238 wl_4 vdd gnd cell_6t
Xbit_r5_c238 bl_238 br_238 wl_5 vdd gnd cell_6t
Xbit_r6_c238 bl_238 br_238 wl_6 vdd gnd cell_6t
Xbit_r7_c238 bl_238 br_238 wl_7 vdd gnd cell_6t
Xbit_r8_c238 bl_238 br_238 wl_8 vdd gnd cell_6t
Xbit_r9_c238 bl_238 br_238 wl_9 vdd gnd cell_6t
Xbit_r10_c238 bl_238 br_238 wl_10 vdd gnd cell_6t
Xbit_r11_c238 bl_238 br_238 wl_11 vdd gnd cell_6t
Xbit_r12_c238 bl_238 br_238 wl_12 vdd gnd cell_6t
Xbit_r13_c238 bl_238 br_238 wl_13 vdd gnd cell_6t
Xbit_r14_c238 bl_238 br_238 wl_14 vdd gnd cell_6t
Xbit_r15_c238 bl_238 br_238 wl_15 vdd gnd cell_6t
Xbit_r16_c238 bl_238 br_238 wl_16 vdd gnd cell_6t
Xbit_r17_c238 bl_238 br_238 wl_17 vdd gnd cell_6t
Xbit_r18_c238 bl_238 br_238 wl_18 vdd gnd cell_6t
Xbit_r19_c238 bl_238 br_238 wl_19 vdd gnd cell_6t
Xbit_r20_c238 bl_238 br_238 wl_20 vdd gnd cell_6t
Xbit_r21_c238 bl_238 br_238 wl_21 vdd gnd cell_6t
Xbit_r22_c238 bl_238 br_238 wl_22 vdd gnd cell_6t
Xbit_r23_c238 bl_238 br_238 wl_23 vdd gnd cell_6t
Xbit_r24_c238 bl_238 br_238 wl_24 vdd gnd cell_6t
Xbit_r25_c238 bl_238 br_238 wl_25 vdd gnd cell_6t
Xbit_r26_c238 bl_238 br_238 wl_26 vdd gnd cell_6t
Xbit_r27_c238 bl_238 br_238 wl_27 vdd gnd cell_6t
Xbit_r28_c238 bl_238 br_238 wl_28 vdd gnd cell_6t
Xbit_r29_c238 bl_238 br_238 wl_29 vdd gnd cell_6t
Xbit_r30_c238 bl_238 br_238 wl_30 vdd gnd cell_6t
Xbit_r31_c238 bl_238 br_238 wl_31 vdd gnd cell_6t
Xbit_r32_c238 bl_238 br_238 wl_32 vdd gnd cell_6t
Xbit_r33_c238 bl_238 br_238 wl_33 vdd gnd cell_6t
Xbit_r34_c238 bl_238 br_238 wl_34 vdd gnd cell_6t
Xbit_r35_c238 bl_238 br_238 wl_35 vdd gnd cell_6t
Xbit_r36_c238 bl_238 br_238 wl_36 vdd gnd cell_6t
Xbit_r37_c238 bl_238 br_238 wl_37 vdd gnd cell_6t
Xbit_r38_c238 bl_238 br_238 wl_38 vdd gnd cell_6t
Xbit_r39_c238 bl_238 br_238 wl_39 vdd gnd cell_6t
Xbit_r40_c238 bl_238 br_238 wl_40 vdd gnd cell_6t
Xbit_r41_c238 bl_238 br_238 wl_41 vdd gnd cell_6t
Xbit_r42_c238 bl_238 br_238 wl_42 vdd gnd cell_6t
Xbit_r43_c238 bl_238 br_238 wl_43 vdd gnd cell_6t
Xbit_r44_c238 bl_238 br_238 wl_44 vdd gnd cell_6t
Xbit_r45_c238 bl_238 br_238 wl_45 vdd gnd cell_6t
Xbit_r46_c238 bl_238 br_238 wl_46 vdd gnd cell_6t
Xbit_r47_c238 bl_238 br_238 wl_47 vdd gnd cell_6t
Xbit_r48_c238 bl_238 br_238 wl_48 vdd gnd cell_6t
Xbit_r49_c238 bl_238 br_238 wl_49 vdd gnd cell_6t
Xbit_r50_c238 bl_238 br_238 wl_50 vdd gnd cell_6t
Xbit_r51_c238 bl_238 br_238 wl_51 vdd gnd cell_6t
Xbit_r52_c238 bl_238 br_238 wl_52 vdd gnd cell_6t
Xbit_r53_c238 bl_238 br_238 wl_53 vdd gnd cell_6t
Xbit_r54_c238 bl_238 br_238 wl_54 vdd gnd cell_6t
Xbit_r55_c238 bl_238 br_238 wl_55 vdd gnd cell_6t
Xbit_r56_c238 bl_238 br_238 wl_56 vdd gnd cell_6t
Xbit_r57_c238 bl_238 br_238 wl_57 vdd gnd cell_6t
Xbit_r58_c238 bl_238 br_238 wl_58 vdd gnd cell_6t
Xbit_r59_c238 bl_238 br_238 wl_59 vdd gnd cell_6t
Xbit_r60_c238 bl_238 br_238 wl_60 vdd gnd cell_6t
Xbit_r61_c238 bl_238 br_238 wl_61 vdd gnd cell_6t
Xbit_r62_c238 bl_238 br_238 wl_62 vdd gnd cell_6t
Xbit_r63_c238 bl_238 br_238 wl_63 vdd gnd cell_6t
Xbit_r64_c238 bl_238 br_238 wl_64 vdd gnd cell_6t
Xbit_r65_c238 bl_238 br_238 wl_65 vdd gnd cell_6t
Xbit_r66_c238 bl_238 br_238 wl_66 vdd gnd cell_6t
Xbit_r67_c238 bl_238 br_238 wl_67 vdd gnd cell_6t
Xbit_r68_c238 bl_238 br_238 wl_68 vdd gnd cell_6t
Xbit_r69_c238 bl_238 br_238 wl_69 vdd gnd cell_6t
Xbit_r70_c238 bl_238 br_238 wl_70 vdd gnd cell_6t
Xbit_r71_c238 bl_238 br_238 wl_71 vdd gnd cell_6t
Xbit_r72_c238 bl_238 br_238 wl_72 vdd gnd cell_6t
Xbit_r73_c238 bl_238 br_238 wl_73 vdd gnd cell_6t
Xbit_r74_c238 bl_238 br_238 wl_74 vdd gnd cell_6t
Xbit_r75_c238 bl_238 br_238 wl_75 vdd gnd cell_6t
Xbit_r76_c238 bl_238 br_238 wl_76 vdd gnd cell_6t
Xbit_r77_c238 bl_238 br_238 wl_77 vdd gnd cell_6t
Xbit_r78_c238 bl_238 br_238 wl_78 vdd gnd cell_6t
Xbit_r79_c238 bl_238 br_238 wl_79 vdd gnd cell_6t
Xbit_r80_c238 bl_238 br_238 wl_80 vdd gnd cell_6t
Xbit_r81_c238 bl_238 br_238 wl_81 vdd gnd cell_6t
Xbit_r82_c238 bl_238 br_238 wl_82 vdd gnd cell_6t
Xbit_r83_c238 bl_238 br_238 wl_83 vdd gnd cell_6t
Xbit_r84_c238 bl_238 br_238 wl_84 vdd gnd cell_6t
Xbit_r85_c238 bl_238 br_238 wl_85 vdd gnd cell_6t
Xbit_r86_c238 bl_238 br_238 wl_86 vdd gnd cell_6t
Xbit_r87_c238 bl_238 br_238 wl_87 vdd gnd cell_6t
Xbit_r88_c238 bl_238 br_238 wl_88 vdd gnd cell_6t
Xbit_r89_c238 bl_238 br_238 wl_89 vdd gnd cell_6t
Xbit_r90_c238 bl_238 br_238 wl_90 vdd gnd cell_6t
Xbit_r91_c238 bl_238 br_238 wl_91 vdd gnd cell_6t
Xbit_r92_c238 bl_238 br_238 wl_92 vdd gnd cell_6t
Xbit_r93_c238 bl_238 br_238 wl_93 vdd gnd cell_6t
Xbit_r94_c238 bl_238 br_238 wl_94 vdd gnd cell_6t
Xbit_r95_c238 bl_238 br_238 wl_95 vdd gnd cell_6t
Xbit_r96_c238 bl_238 br_238 wl_96 vdd gnd cell_6t
Xbit_r97_c238 bl_238 br_238 wl_97 vdd gnd cell_6t
Xbit_r98_c238 bl_238 br_238 wl_98 vdd gnd cell_6t
Xbit_r99_c238 bl_238 br_238 wl_99 vdd gnd cell_6t
Xbit_r100_c238 bl_238 br_238 wl_100 vdd gnd cell_6t
Xbit_r101_c238 bl_238 br_238 wl_101 vdd gnd cell_6t
Xbit_r102_c238 bl_238 br_238 wl_102 vdd gnd cell_6t
Xbit_r103_c238 bl_238 br_238 wl_103 vdd gnd cell_6t
Xbit_r104_c238 bl_238 br_238 wl_104 vdd gnd cell_6t
Xbit_r105_c238 bl_238 br_238 wl_105 vdd gnd cell_6t
Xbit_r106_c238 bl_238 br_238 wl_106 vdd gnd cell_6t
Xbit_r107_c238 bl_238 br_238 wl_107 vdd gnd cell_6t
Xbit_r108_c238 bl_238 br_238 wl_108 vdd gnd cell_6t
Xbit_r109_c238 bl_238 br_238 wl_109 vdd gnd cell_6t
Xbit_r110_c238 bl_238 br_238 wl_110 vdd gnd cell_6t
Xbit_r111_c238 bl_238 br_238 wl_111 vdd gnd cell_6t
Xbit_r112_c238 bl_238 br_238 wl_112 vdd gnd cell_6t
Xbit_r113_c238 bl_238 br_238 wl_113 vdd gnd cell_6t
Xbit_r114_c238 bl_238 br_238 wl_114 vdd gnd cell_6t
Xbit_r115_c238 bl_238 br_238 wl_115 vdd gnd cell_6t
Xbit_r116_c238 bl_238 br_238 wl_116 vdd gnd cell_6t
Xbit_r117_c238 bl_238 br_238 wl_117 vdd gnd cell_6t
Xbit_r118_c238 bl_238 br_238 wl_118 vdd gnd cell_6t
Xbit_r119_c238 bl_238 br_238 wl_119 vdd gnd cell_6t
Xbit_r120_c238 bl_238 br_238 wl_120 vdd gnd cell_6t
Xbit_r121_c238 bl_238 br_238 wl_121 vdd gnd cell_6t
Xbit_r122_c238 bl_238 br_238 wl_122 vdd gnd cell_6t
Xbit_r123_c238 bl_238 br_238 wl_123 vdd gnd cell_6t
Xbit_r124_c238 bl_238 br_238 wl_124 vdd gnd cell_6t
Xbit_r125_c238 bl_238 br_238 wl_125 vdd gnd cell_6t
Xbit_r126_c238 bl_238 br_238 wl_126 vdd gnd cell_6t
Xbit_r127_c238 bl_238 br_238 wl_127 vdd gnd cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd cell_6t
Xbit_r1_c239 bl_239 br_239 wl_1 vdd gnd cell_6t
Xbit_r2_c239 bl_239 br_239 wl_2 vdd gnd cell_6t
Xbit_r3_c239 bl_239 br_239 wl_3 vdd gnd cell_6t
Xbit_r4_c239 bl_239 br_239 wl_4 vdd gnd cell_6t
Xbit_r5_c239 bl_239 br_239 wl_5 vdd gnd cell_6t
Xbit_r6_c239 bl_239 br_239 wl_6 vdd gnd cell_6t
Xbit_r7_c239 bl_239 br_239 wl_7 vdd gnd cell_6t
Xbit_r8_c239 bl_239 br_239 wl_8 vdd gnd cell_6t
Xbit_r9_c239 bl_239 br_239 wl_9 vdd gnd cell_6t
Xbit_r10_c239 bl_239 br_239 wl_10 vdd gnd cell_6t
Xbit_r11_c239 bl_239 br_239 wl_11 vdd gnd cell_6t
Xbit_r12_c239 bl_239 br_239 wl_12 vdd gnd cell_6t
Xbit_r13_c239 bl_239 br_239 wl_13 vdd gnd cell_6t
Xbit_r14_c239 bl_239 br_239 wl_14 vdd gnd cell_6t
Xbit_r15_c239 bl_239 br_239 wl_15 vdd gnd cell_6t
Xbit_r16_c239 bl_239 br_239 wl_16 vdd gnd cell_6t
Xbit_r17_c239 bl_239 br_239 wl_17 vdd gnd cell_6t
Xbit_r18_c239 bl_239 br_239 wl_18 vdd gnd cell_6t
Xbit_r19_c239 bl_239 br_239 wl_19 vdd gnd cell_6t
Xbit_r20_c239 bl_239 br_239 wl_20 vdd gnd cell_6t
Xbit_r21_c239 bl_239 br_239 wl_21 vdd gnd cell_6t
Xbit_r22_c239 bl_239 br_239 wl_22 vdd gnd cell_6t
Xbit_r23_c239 bl_239 br_239 wl_23 vdd gnd cell_6t
Xbit_r24_c239 bl_239 br_239 wl_24 vdd gnd cell_6t
Xbit_r25_c239 bl_239 br_239 wl_25 vdd gnd cell_6t
Xbit_r26_c239 bl_239 br_239 wl_26 vdd gnd cell_6t
Xbit_r27_c239 bl_239 br_239 wl_27 vdd gnd cell_6t
Xbit_r28_c239 bl_239 br_239 wl_28 vdd gnd cell_6t
Xbit_r29_c239 bl_239 br_239 wl_29 vdd gnd cell_6t
Xbit_r30_c239 bl_239 br_239 wl_30 vdd gnd cell_6t
Xbit_r31_c239 bl_239 br_239 wl_31 vdd gnd cell_6t
Xbit_r32_c239 bl_239 br_239 wl_32 vdd gnd cell_6t
Xbit_r33_c239 bl_239 br_239 wl_33 vdd gnd cell_6t
Xbit_r34_c239 bl_239 br_239 wl_34 vdd gnd cell_6t
Xbit_r35_c239 bl_239 br_239 wl_35 vdd gnd cell_6t
Xbit_r36_c239 bl_239 br_239 wl_36 vdd gnd cell_6t
Xbit_r37_c239 bl_239 br_239 wl_37 vdd gnd cell_6t
Xbit_r38_c239 bl_239 br_239 wl_38 vdd gnd cell_6t
Xbit_r39_c239 bl_239 br_239 wl_39 vdd gnd cell_6t
Xbit_r40_c239 bl_239 br_239 wl_40 vdd gnd cell_6t
Xbit_r41_c239 bl_239 br_239 wl_41 vdd gnd cell_6t
Xbit_r42_c239 bl_239 br_239 wl_42 vdd gnd cell_6t
Xbit_r43_c239 bl_239 br_239 wl_43 vdd gnd cell_6t
Xbit_r44_c239 bl_239 br_239 wl_44 vdd gnd cell_6t
Xbit_r45_c239 bl_239 br_239 wl_45 vdd gnd cell_6t
Xbit_r46_c239 bl_239 br_239 wl_46 vdd gnd cell_6t
Xbit_r47_c239 bl_239 br_239 wl_47 vdd gnd cell_6t
Xbit_r48_c239 bl_239 br_239 wl_48 vdd gnd cell_6t
Xbit_r49_c239 bl_239 br_239 wl_49 vdd gnd cell_6t
Xbit_r50_c239 bl_239 br_239 wl_50 vdd gnd cell_6t
Xbit_r51_c239 bl_239 br_239 wl_51 vdd gnd cell_6t
Xbit_r52_c239 bl_239 br_239 wl_52 vdd gnd cell_6t
Xbit_r53_c239 bl_239 br_239 wl_53 vdd gnd cell_6t
Xbit_r54_c239 bl_239 br_239 wl_54 vdd gnd cell_6t
Xbit_r55_c239 bl_239 br_239 wl_55 vdd gnd cell_6t
Xbit_r56_c239 bl_239 br_239 wl_56 vdd gnd cell_6t
Xbit_r57_c239 bl_239 br_239 wl_57 vdd gnd cell_6t
Xbit_r58_c239 bl_239 br_239 wl_58 vdd gnd cell_6t
Xbit_r59_c239 bl_239 br_239 wl_59 vdd gnd cell_6t
Xbit_r60_c239 bl_239 br_239 wl_60 vdd gnd cell_6t
Xbit_r61_c239 bl_239 br_239 wl_61 vdd gnd cell_6t
Xbit_r62_c239 bl_239 br_239 wl_62 vdd gnd cell_6t
Xbit_r63_c239 bl_239 br_239 wl_63 vdd gnd cell_6t
Xbit_r64_c239 bl_239 br_239 wl_64 vdd gnd cell_6t
Xbit_r65_c239 bl_239 br_239 wl_65 vdd gnd cell_6t
Xbit_r66_c239 bl_239 br_239 wl_66 vdd gnd cell_6t
Xbit_r67_c239 bl_239 br_239 wl_67 vdd gnd cell_6t
Xbit_r68_c239 bl_239 br_239 wl_68 vdd gnd cell_6t
Xbit_r69_c239 bl_239 br_239 wl_69 vdd gnd cell_6t
Xbit_r70_c239 bl_239 br_239 wl_70 vdd gnd cell_6t
Xbit_r71_c239 bl_239 br_239 wl_71 vdd gnd cell_6t
Xbit_r72_c239 bl_239 br_239 wl_72 vdd gnd cell_6t
Xbit_r73_c239 bl_239 br_239 wl_73 vdd gnd cell_6t
Xbit_r74_c239 bl_239 br_239 wl_74 vdd gnd cell_6t
Xbit_r75_c239 bl_239 br_239 wl_75 vdd gnd cell_6t
Xbit_r76_c239 bl_239 br_239 wl_76 vdd gnd cell_6t
Xbit_r77_c239 bl_239 br_239 wl_77 vdd gnd cell_6t
Xbit_r78_c239 bl_239 br_239 wl_78 vdd gnd cell_6t
Xbit_r79_c239 bl_239 br_239 wl_79 vdd gnd cell_6t
Xbit_r80_c239 bl_239 br_239 wl_80 vdd gnd cell_6t
Xbit_r81_c239 bl_239 br_239 wl_81 vdd gnd cell_6t
Xbit_r82_c239 bl_239 br_239 wl_82 vdd gnd cell_6t
Xbit_r83_c239 bl_239 br_239 wl_83 vdd gnd cell_6t
Xbit_r84_c239 bl_239 br_239 wl_84 vdd gnd cell_6t
Xbit_r85_c239 bl_239 br_239 wl_85 vdd gnd cell_6t
Xbit_r86_c239 bl_239 br_239 wl_86 vdd gnd cell_6t
Xbit_r87_c239 bl_239 br_239 wl_87 vdd gnd cell_6t
Xbit_r88_c239 bl_239 br_239 wl_88 vdd gnd cell_6t
Xbit_r89_c239 bl_239 br_239 wl_89 vdd gnd cell_6t
Xbit_r90_c239 bl_239 br_239 wl_90 vdd gnd cell_6t
Xbit_r91_c239 bl_239 br_239 wl_91 vdd gnd cell_6t
Xbit_r92_c239 bl_239 br_239 wl_92 vdd gnd cell_6t
Xbit_r93_c239 bl_239 br_239 wl_93 vdd gnd cell_6t
Xbit_r94_c239 bl_239 br_239 wl_94 vdd gnd cell_6t
Xbit_r95_c239 bl_239 br_239 wl_95 vdd gnd cell_6t
Xbit_r96_c239 bl_239 br_239 wl_96 vdd gnd cell_6t
Xbit_r97_c239 bl_239 br_239 wl_97 vdd gnd cell_6t
Xbit_r98_c239 bl_239 br_239 wl_98 vdd gnd cell_6t
Xbit_r99_c239 bl_239 br_239 wl_99 vdd gnd cell_6t
Xbit_r100_c239 bl_239 br_239 wl_100 vdd gnd cell_6t
Xbit_r101_c239 bl_239 br_239 wl_101 vdd gnd cell_6t
Xbit_r102_c239 bl_239 br_239 wl_102 vdd gnd cell_6t
Xbit_r103_c239 bl_239 br_239 wl_103 vdd gnd cell_6t
Xbit_r104_c239 bl_239 br_239 wl_104 vdd gnd cell_6t
Xbit_r105_c239 bl_239 br_239 wl_105 vdd gnd cell_6t
Xbit_r106_c239 bl_239 br_239 wl_106 vdd gnd cell_6t
Xbit_r107_c239 bl_239 br_239 wl_107 vdd gnd cell_6t
Xbit_r108_c239 bl_239 br_239 wl_108 vdd gnd cell_6t
Xbit_r109_c239 bl_239 br_239 wl_109 vdd gnd cell_6t
Xbit_r110_c239 bl_239 br_239 wl_110 vdd gnd cell_6t
Xbit_r111_c239 bl_239 br_239 wl_111 vdd gnd cell_6t
Xbit_r112_c239 bl_239 br_239 wl_112 vdd gnd cell_6t
Xbit_r113_c239 bl_239 br_239 wl_113 vdd gnd cell_6t
Xbit_r114_c239 bl_239 br_239 wl_114 vdd gnd cell_6t
Xbit_r115_c239 bl_239 br_239 wl_115 vdd gnd cell_6t
Xbit_r116_c239 bl_239 br_239 wl_116 vdd gnd cell_6t
Xbit_r117_c239 bl_239 br_239 wl_117 vdd gnd cell_6t
Xbit_r118_c239 bl_239 br_239 wl_118 vdd gnd cell_6t
Xbit_r119_c239 bl_239 br_239 wl_119 vdd gnd cell_6t
Xbit_r120_c239 bl_239 br_239 wl_120 vdd gnd cell_6t
Xbit_r121_c239 bl_239 br_239 wl_121 vdd gnd cell_6t
Xbit_r122_c239 bl_239 br_239 wl_122 vdd gnd cell_6t
Xbit_r123_c239 bl_239 br_239 wl_123 vdd gnd cell_6t
Xbit_r124_c239 bl_239 br_239 wl_124 vdd gnd cell_6t
Xbit_r125_c239 bl_239 br_239 wl_125 vdd gnd cell_6t
Xbit_r126_c239 bl_239 br_239 wl_126 vdd gnd cell_6t
Xbit_r127_c239 bl_239 br_239 wl_127 vdd gnd cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd cell_6t
Xbit_r1_c240 bl_240 br_240 wl_1 vdd gnd cell_6t
Xbit_r2_c240 bl_240 br_240 wl_2 vdd gnd cell_6t
Xbit_r3_c240 bl_240 br_240 wl_3 vdd gnd cell_6t
Xbit_r4_c240 bl_240 br_240 wl_4 vdd gnd cell_6t
Xbit_r5_c240 bl_240 br_240 wl_5 vdd gnd cell_6t
Xbit_r6_c240 bl_240 br_240 wl_6 vdd gnd cell_6t
Xbit_r7_c240 bl_240 br_240 wl_7 vdd gnd cell_6t
Xbit_r8_c240 bl_240 br_240 wl_8 vdd gnd cell_6t
Xbit_r9_c240 bl_240 br_240 wl_9 vdd gnd cell_6t
Xbit_r10_c240 bl_240 br_240 wl_10 vdd gnd cell_6t
Xbit_r11_c240 bl_240 br_240 wl_11 vdd gnd cell_6t
Xbit_r12_c240 bl_240 br_240 wl_12 vdd gnd cell_6t
Xbit_r13_c240 bl_240 br_240 wl_13 vdd gnd cell_6t
Xbit_r14_c240 bl_240 br_240 wl_14 vdd gnd cell_6t
Xbit_r15_c240 bl_240 br_240 wl_15 vdd gnd cell_6t
Xbit_r16_c240 bl_240 br_240 wl_16 vdd gnd cell_6t
Xbit_r17_c240 bl_240 br_240 wl_17 vdd gnd cell_6t
Xbit_r18_c240 bl_240 br_240 wl_18 vdd gnd cell_6t
Xbit_r19_c240 bl_240 br_240 wl_19 vdd gnd cell_6t
Xbit_r20_c240 bl_240 br_240 wl_20 vdd gnd cell_6t
Xbit_r21_c240 bl_240 br_240 wl_21 vdd gnd cell_6t
Xbit_r22_c240 bl_240 br_240 wl_22 vdd gnd cell_6t
Xbit_r23_c240 bl_240 br_240 wl_23 vdd gnd cell_6t
Xbit_r24_c240 bl_240 br_240 wl_24 vdd gnd cell_6t
Xbit_r25_c240 bl_240 br_240 wl_25 vdd gnd cell_6t
Xbit_r26_c240 bl_240 br_240 wl_26 vdd gnd cell_6t
Xbit_r27_c240 bl_240 br_240 wl_27 vdd gnd cell_6t
Xbit_r28_c240 bl_240 br_240 wl_28 vdd gnd cell_6t
Xbit_r29_c240 bl_240 br_240 wl_29 vdd gnd cell_6t
Xbit_r30_c240 bl_240 br_240 wl_30 vdd gnd cell_6t
Xbit_r31_c240 bl_240 br_240 wl_31 vdd gnd cell_6t
Xbit_r32_c240 bl_240 br_240 wl_32 vdd gnd cell_6t
Xbit_r33_c240 bl_240 br_240 wl_33 vdd gnd cell_6t
Xbit_r34_c240 bl_240 br_240 wl_34 vdd gnd cell_6t
Xbit_r35_c240 bl_240 br_240 wl_35 vdd gnd cell_6t
Xbit_r36_c240 bl_240 br_240 wl_36 vdd gnd cell_6t
Xbit_r37_c240 bl_240 br_240 wl_37 vdd gnd cell_6t
Xbit_r38_c240 bl_240 br_240 wl_38 vdd gnd cell_6t
Xbit_r39_c240 bl_240 br_240 wl_39 vdd gnd cell_6t
Xbit_r40_c240 bl_240 br_240 wl_40 vdd gnd cell_6t
Xbit_r41_c240 bl_240 br_240 wl_41 vdd gnd cell_6t
Xbit_r42_c240 bl_240 br_240 wl_42 vdd gnd cell_6t
Xbit_r43_c240 bl_240 br_240 wl_43 vdd gnd cell_6t
Xbit_r44_c240 bl_240 br_240 wl_44 vdd gnd cell_6t
Xbit_r45_c240 bl_240 br_240 wl_45 vdd gnd cell_6t
Xbit_r46_c240 bl_240 br_240 wl_46 vdd gnd cell_6t
Xbit_r47_c240 bl_240 br_240 wl_47 vdd gnd cell_6t
Xbit_r48_c240 bl_240 br_240 wl_48 vdd gnd cell_6t
Xbit_r49_c240 bl_240 br_240 wl_49 vdd gnd cell_6t
Xbit_r50_c240 bl_240 br_240 wl_50 vdd gnd cell_6t
Xbit_r51_c240 bl_240 br_240 wl_51 vdd gnd cell_6t
Xbit_r52_c240 bl_240 br_240 wl_52 vdd gnd cell_6t
Xbit_r53_c240 bl_240 br_240 wl_53 vdd gnd cell_6t
Xbit_r54_c240 bl_240 br_240 wl_54 vdd gnd cell_6t
Xbit_r55_c240 bl_240 br_240 wl_55 vdd gnd cell_6t
Xbit_r56_c240 bl_240 br_240 wl_56 vdd gnd cell_6t
Xbit_r57_c240 bl_240 br_240 wl_57 vdd gnd cell_6t
Xbit_r58_c240 bl_240 br_240 wl_58 vdd gnd cell_6t
Xbit_r59_c240 bl_240 br_240 wl_59 vdd gnd cell_6t
Xbit_r60_c240 bl_240 br_240 wl_60 vdd gnd cell_6t
Xbit_r61_c240 bl_240 br_240 wl_61 vdd gnd cell_6t
Xbit_r62_c240 bl_240 br_240 wl_62 vdd gnd cell_6t
Xbit_r63_c240 bl_240 br_240 wl_63 vdd gnd cell_6t
Xbit_r64_c240 bl_240 br_240 wl_64 vdd gnd cell_6t
Xbit_r65_c240 bl_240 br_240 wl_65 vdd gnd cell_6t
Xbit_r66_c240 bl_240 br_240 wl_66 vdd gnd cell_6t
Xbit_r67_c240 bl_240 br_240 wl_67 vdd gnd cell_6t
Xbit_r68_c240 bl_240 br_240 wl_68 vdd gnd cell_6t
Xbit_r69_c240 bl_240 br_240 wl_69 vdd gnd cell_6t
Xbit_r70_c240 bl_240 br_240 wl_70 vdd gnd cell_6t
Xbit_r71_c240 bl_240 br_240 wl_71 vdd gnd cell_6t
Xbit_r72_c240 bl_240 br_240 wl_72 vdd gnd cell_6t
Xbit_r73_c240 bl_240 br_240 wl_73 vdd gnd cell_6t
Xbit_r74_c240 bl_240 br_240 wl_74 vdd gnd cell_6t
Xbit_r75_c240 bl_240 br_240 wl_75 vdd gnd cell_6t
Xbit_r76_c240 bl_240 br_240 wl_76 vdd gnd cell_6t
Xbit_r77_c240 bl_240 br_240 wl_77 vdd gnd cell_6t
Xbit_r78_c240 bl_240 br_240 wl_78 vdd gnd cell_6t
Xbit_r79_c240 bl_240 br_240 wl_79 vdd gnd cell_6t
Xbit_r80_c240 bl_240 br_240 wl_80 vdd gnd cell_6t
Xbit_r81_c240 bl_240 br_240 wl_81 vdd gnd cell_6t
Xbit_r82_c240 bl_240 br_240 wl_82 vdd gnd cell_6t
Xbit_r83_c240 bl_240 br_240 wl_83 vdd gnd cell_6t
Xbit_r84_c240 bl_240 br_240 wl_84 vdd gnd cell_6t
Xbit_r85_c240 bl_240 br_240 wl_85 vdd gnd cell_6t
Xbit_r86_c240 bl_240 br_240 wl_86 vdd gnd cell_6t
Xbit_r87_c240 bl_240 br_240 wl_87 vdd gnd cell_6t
Xbit_r88_c240 bl_240 br_240 wl_88 vdd gnd cell_6t
Xbit_r89_c240 bl_240 br_240 wl_89 vdd gnd cell_6t
Xbit_r90_c240 bl_240 br_240 wl_90 vdd gnd cell_6t
Xbit_r91_c240 bl_240 br_240 wl_91 vdd gnd cell_6t
Xbit_r92_c240 bl_240 br_240 wl_92 vdd gnd cell_6t
Xbit_r93_c240 bl_240 br_240 wl_93 vdd gnd cell_6t
Xbit_r94_c240 bl_240 br_240 wl_94 vdd gnd cell_6t
Xbit_r95_c240 bl_240 br_240 wl_95 vdd gnd cell_6t
Xbit_r96_c240 bl_240 br_240 wl_96 vdd gnd cell_6t
Xbit_r97_c240 bl_240 br_240 wl_97 vdd gnd cell_6t
Xbit_r98_c240 bl_240 br_240 wl_98 vdd gnd cell_6t
Xbit_r99_c240 bl_240 br_240 wl_99 vdd gnd cell_6t
Xbit_r100_c240 bl_240 br_240 wl_100 vdd gnd cell_6t
Xbit_r101_c240 bl_240 br_240 wl_101 vdd gnd cell_6t
Xbit_r102_c240 bl_240 br_240 wl_102 vdd gnd cell_6t
Xbit_r103_c240 bl_240 br_240 wl_103 vdd gnd cell_6t
Xbit_r104_c240 bl_240 br_240 wl_104 vdd gnd cell_6t
Xbit_r105_c240 bl_240 br_240 wl_105 vdd gnd cell_6t
Xbit_r106_c240 bl_240 br_240 wl_106 vdd gnd cell_6t
Xbit_r107_c240 bl_240 br_240 wl_107 vdd gnd cell_6t
Xbit_r108_c240 bl_240 br_240 wl_108 vdd gnd cell_6t
Xbit_r109_c240 bl_240 br_240 wl_109 vdd gnd cell_6t
Xbit_r110_c240 bl_240 br_240 wl_110 vdd gnd cell_6t
Xbit_r111_c240 bl_240 br_240 wl_111 vdd gnd cell_6t
Xbit_r112_c240 bl_240 br_240 wl_112 vdd gnd cell_6t
Xbit_r113_c240 bl_240 br_240 wl_113 vdd gnd cell_6t
Xbit_r114_c240 bl_240 br_240 wl_114 vdd gnd cell_6t
Xbit_r115_c240 bl_240 br_240 wl_115 vdd gnd cell_6t
Xbit_r116_c240 bl_240 br_240 wl_116 vdd gnd cell_6t
Xbit_r117_c240 bl_240 br_240 wl_117 vdd gnd cell_6t
Xbit_r118_c240 bl_240 br_240 wl_118 vdd gnd cell_6t
Xbit_r119_c240 bl_240 br_240 wl_119 vdd gnd cell_6t
Xbit_r120_c240 bl_240 br_240 wl_120 vdd gnd cell_6t
Xbit_r121_c240 bl_240 br_240 wl_121 vdd gnd cell_6t
Xbit_r122_c240 bl_240 br_240 wl_122 vdd gnd cell_6t
Xbit_r123_c240 bl_240 br_240 wl_123 vdd gnd cell_6t
Xbit_r124_c240 bl_240 br_240 wl_124 vdd gnd cell_6t
Xbit_r125_c240 bl_240 br_240 wl_125 vdd gnd cell_6t
Xbit_r126_c240 bl_240 br_240 wl_126 vdd gnd cell_6t
Xbit_r127_c240 bl_240 br_240 wl_127 vdd gnd cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd cell_6t
Xbit_r1_c241 bl_241 br_241 wl_1 vdd gnd cell_6t
Xbit_r2_c241 bl_241 br_241 wl_2 vdd gnd cell_6t
Xbit_r3_c241 bl_241 br_241 wl_3 vdd gnd cell_6t
Xbit_r4_c241 bl_241 br_241 wl_4 vdd gnd cell_6t
Xbit_r5_c241 bl_241 br_241 wl_5 vdd gnd cell_6t
Xbit_r6_c241 bl_241 br_241 wl_6 vdd gnd cell_6t
Xbit_r7_c241 bl_241 br_241 wl_7 vdd gnd cell_6t
Xbit_r8_c241 bl_241 br_241 wl_8 vdd gnd cell_6t
Xbit_r9_c241 bl_241 br_241 wl_9 vdd gnd cell_6t
Xbit_r10_c241 bl_241 br_241 wl_10 vdd gnd cell_6t
Xbit_r11_c241 bl_241 br_241 wl_11 vdd gnd cell_6t
Xbit_r12_c241 bl_241 br_241 wl_12 vdd gnd cell_6t
Xbit_r13_c241 bl_241 br_241 wl_13 vdd gnd cell_6t
Xbit_r14_c241 bl_241 br_241 wl_14 vdd gnd cell_6t
Xbit_r15_c241 bl_241 br_241 wl_15 vdd gnd cell_6t
Xbit_r16_c241 bl_241 br_241 wl_16 vdd gnd cell_6t
Xbit_r17_c241 bl_241 br_241 wl_17 vdd gnd cell_6t
Xbit_r18_c241 bl_241 br_241 wl_18 vdd gnd cell_6t
Xbit_r19_c241 bl_241 br_241 wl_19 vdd gnd cell_6t
Xbit_r20_c241 bl_241 br_241 wl_20 vdd gnd cell_6t
Xbit_r21_c241 bl_241 br_241 wl_21 vdd gnd cell_6t
Xbit_r22_c241 bl_241 br_241 wl_22 vdd gnd cell_6t
Xbit_r23_c241 bl_241 br_241 wl_23 vdd gnd cell_6t
Xbit_r24_c241 bl_241 br_241 wl_24 vdd gnd cell_6t
Xbit_r25_c241 bl_241 br_241 wl_25 vdd gnd cell_6t
Xbit_r26_c241 bl_241 br_241 wl_26 vdd gnd cell_6t
Xbit_r27_c241 bl_241 br_241 wl_27 vdd gnd cell_6t
Xbit_r28_c241 bl_241 br_241 wl_28 vdd gnd cell_6t
Xbit_r29_c241 bl_241 br_241 wl_29 vdd gnd cell_6t
Xbit_r30_c241 bl_241 br_241 wl_30 vdd gnd cell_6t
Xbit_r31_c241 bl_241 br_241 wl_31 vdd gnd cell_6t
Xbit_r32_c241 bl_241 br_241 wl_32 vdd gnd cell_6t
Xbit_r33_c241 bl_241 br_241 wl_33 vdd gnd cell_6t
Xbit_r34_c241 bl_241 br_241 wl_34 vdd gnd cell_6t
Xbit_r35_c241 bl_241 br_241 wl_35 vdd gnd cell_6t
Xbit_r36_c241 bl_241 br_241 wl_36 vdd gnd cell_6t
Xbit_r37_c241 bl_241 br_241 wl_37 vdd gnd cell_6t
Xbit_r38_c241 bl_241 br_241 wl_38 vdd gnd cell_6t
Xbit_r39_c241 bl_241 br_241 wl_39 vdd gnd cell_6t
Xbit_r40_c241 bl_241 br_241 wl_40 vdd gnd cell_6t
Xbit_r41_c241 bl_241 br_241 wl_41 vdd gnd cell_6t
Xbit_r42_c241 bl_241 br_241 wl_42 vdd gnd cell_6t
Xbit_r43_c241 bl_241 br_241 wl_43 vdd gnd cell_6t
Xbit_r44_c241 bl_241 br_241 wl_44 vdd gnd cell_6t
Xbit_r45_c241 bl_241 br_241 wl_45 vdd gnd cell_6t
Xbit_r46_c241 bl_241 br_241 wl_46 vdd gnd cell_6t
Xbit_r47_c241 bl_241 br_241 wl_47 vdd gnd cell_6t
Xbit_r48_c241 bl_241 br_241 wl_48 vdd gnd cell_6t
Xbit_r49_c241 bl_241 br_241 wl_49 vdd gnd cell_6t
Xbit_r50_c241 bl_241 br_241 wl_50 vdd gnd cell_6t
Xbit_r51_c241 bl_241 br_241 wl_51 vdd gnd cell_6t
Xbit_r52_c241 bl_241 br_241 wl_52 vdd gnd cell_6t
Xbit_r53_c241 bl_241 br_241 wl_53 vdd gnd cell_6t
Xbit_r54_c241 bl_241 br_241 wl_54 vdd gnd cell_6t
Xbit_r55_c241 bl_241 br_241 wl_55 vdd gnd cell_6t
Xbit_r56_c241 bl_241 br_241 wl_56 vdd gnd cell_6t
Xbit_r57_c241 bl_241 br_241 wl_57 vdd gnd cell_6t
Xbit_r58_c241 bl_241 br_241 wl_58 vdd gnd cell_6t
Xbit_r59_c241 bl_241 br_241 wl_59 vdd gnd cell_6t
Xbit_r60_c241 bl_241 br_241 wl_60 vdd gnd cell_6t
Xbit_r61_c241 bl_241 br_241 wl_61 vdd gnd cell_6t
Xbit_r62_c241 bl_241 br_241 wl_62 vdd gnd cell_6t
Xbit_r63_c241 bl_241 br_241 wl_63 vdd gnd cell_6t
Xbit_r64_c241 bl_241 br_241 wl_64 vdd gnd cell_6t
Xbit_r65_c241 bl_241 br_241 wl_65 vdd gnd cell_6t
Xbit_r66_c241 bl_241 br_241 wl_66 vdd gnd cell_6t
Xbit_r67_c241 bl_241 br_241 wl_67 vdd gnd cell_6t
Xbit_r68_c241 bl_241 br_241 wl_68 vdd gnd cell_6t
Xbit_r69_c241 bl_241 br_241 wl_69 vdd gnd cell_6t
Xbit_r70_c241 bl_241 br_241 wl_70 vdd gnd cell_6t
Xbit_r71_c241 bl_241 br_241 wl_71 vdd gnd cell_6t
Xbit_r72_c241 bl_241 br_241 wl_72 vdd gnd cell_6t
Xbit_r73_c241 bl_241 br_241 wl_73 vdd gnd cell_6t
Xbit_r74_c241 bl_241 br_241 wl_74 vdd gnd cell_6t
Xbit_r75_c241 bl_241 br_241 wl_75 vdd gnd cell_6t
Xbit_r76_c241 bl_241 br_241 wl_76 vdd gnd cell_6t
Xbit_r77_c241 bl_241 br_241 wl_77 vdd gnd cell_6t
Xbit_r78_c241 bl_241 br_241 wl_78 vdd gnd cell_6t
Xbit_r79_c241 bl_241 br_241 wl_79 vdd gnd cell_6t
Xbit_r80_c241 bl_241 br_241 wl_80 vdd gnd cell_6t
Xbit_r81_c241 bl_241 br_241 wl_81 vdd gnd cell_6t
Xbit_r82_c241 bl_241 br_241 wl_82 vdd gnd cell_6t
Xbit_r83_c241 bl_241 br_241 wl_83 vdd gnd cell_6t
Xbit_r84_c241 bl_241 br_241 wl_84 vdd gnd cell_6t
Xbit_r85_c241 bl_241 br_241 wl_85 vdd gnd cell_6t
Xbit_r86_c241 bl_241 br_241 wl_86 vdd gnd cell_6t
Xbit_r87_c241 bl_241 br_241 wl_87 vdd gnd cell_6t
Xbit_r88_c241 bl_241 br_241 wl_88 vdd gnd cell_6t
Xbit_r89_c241 bl_241 br_241 wl_89 vdd gnd cell_6t
Xbit_r90_c241 bl_241 br_241 wl_90 vdd gnd cell_6t
Xbit_r91_c241 bl_241 br_241 wl_91 vdd gnd cell_6t
Xbit_r92_c241 bl_241 br_241 wl_92 vdd gnd cell_6t
Xbit_r93_c241 bl_241 br_241 wl_93 vdd gnd cell_6t
Xbit_r94_c241 bl_241 br_241 wl_94 vdd gnd cell_6t
Xbit_r95_c241 bl_241 br_241 wl_95 vdd gnd cell_6t
Xbit_r96_c241 bl_241 br_241 wl_96 vdd gnd cell_6t
Xbit_r97_c241 bl_241 br_241 wl_97 vdd gnd cell_6t
Xbit_r98_c241 bl_241 br_241 wl_98 vdd gnd cell_6t
Xbit_r99_c241 bl_241 br_241 wl_99 vdd gnd cell_6t
Xbit_r100_c241 bl_241 br_241 wl_100 vdd gnd cell_6t
Xbit_r101_c241 bl_241 br_241 wl_101 vdd gnd cell_6t
Xbit_r102_c241 bl_241 br_241 wl_102 vdd gnd cell_6t
Xbit_r103_c241 bl_241 br_241 wl_103 vdd gnd cell_6t
Xbit_r104_c241 bl_241 br_241 wl_104 vdd gnd cell_6t
Xbit_r105_c241 bl_241 br_241 wl_105 vdd gnd cell_6t
Xbit_r106_c241 bl_241 br_241 wl_106 vdd gnd cell_6t
Xbit_r107_c241 bl_241 br_241 wl_107 vdd gnd cell_6t
Xbit_r108_c241 bl_241 br_241 wl_108 vdd gnd cell_6t
Xbit_r109_c241 bl_241 br_241 wl_109 vdd gnd cell_6t
Xbit_r110_c241 bl_241 br_241 wl_110 vdd gnd cell_6t
Xbit_r111_c241 bl_241 br_241 wl_111 vdd gnd cell_6t
Xbit_r112_c241 bl_241 br_241 wl_112 vdd gnd cell_6t
Xbit_r113_c241 bl_241 br_241 wl_113 vdd gnd cell_6t
Xbit_r114_c241 bl_241 br_241 wl_114 vdd gnd cell_6t
Xbit_r115_c241 bl_241 br_241 wl_115 vdd gnd cell_6t
Xbit_r116_c241 bl_241 br_241 wl_116 vdd gnd cell_6t
Xbit_r117_c241 bl_241 br_241 wl_117 vdd gnd cell_6t
Xbit_r118_c241 bl_241 br_241 wl_118 vdd gnd cell_6t
Xbit_r119_c241 bl_241 br_241 wl_119 vdd gnd cell_6t
Xbit_r120_c241 bl_241 br_241 wl_120 vdd gnd cell_6t
Xbit_r121_c241 bl_241 br_241 wl_121 vdd gnd cell_6t
Xbit_r122_c241 bl_241 br_241 wl_122 vdd gnd cell_6t
Xbit_r123_c241 bl_241 br_241 wl_123 vdd gnd cell_6t
Xbit_r124_c241 bl_241 br_241 wl_124 vdd gnd cell_6t
Xbit_r125_c241 bl_241 br_241 wl_125 vdd gnd cell_6t
Xbit_r126_c241 bl_241 br_241 wl_126 vdd gnd cell_6t
Xbit_r127_c241 bl_241 br_241 wl_127 vdd gnd cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd cell_6t
Xbit_r1_c242 bl_242 br_242 wl_1 vdd gnd cell_6t
Xbit_r2_c242 bl_242 br_242 wl_2 vdd gnd cell_6t
Xbit_r3_c242 bl_242 br_242 wl_3 vdd gnd cell_6t
Xbit_r4_c242 bl_242 br_242 wl_4 vdd gnd cell_6t
Xbit_r5_c242 bl_242 br_242 wl_5 vdd gnd cell_6t
Xbit_r6_c242 bl_242 br_242 wl_6 vdd gnd cell_6t
Xbit_r7_c242 bl_242 br_242 wl_7 vdd gnd cell_6t
Xbit_r8_c242 bl_242 br_242 wl_8 vdd gnd cell_6t
Xbit_r9_c242 bl_242 br_242 wl_9 vdd gnd cell_6t
Xbit_r10_c242 bl_242 br_242 wl_10 vdd gnd cell_6t
Xbit_r11_c242 bl_242 br_242 wl_11 vdd gnd cell_6t
Xbit_r12_c242 bl_242 br_242 wl_12 vdd gnd cell_6t
Xbit_r13_c242 bl_242 br_242 wl_13 vdd gnd cell_6t
Xbit_r14_c242 bl_242 br_242 wl_14 vdd gnd cell_6t
Xbit_r15_c242 bl_242 br_242 wl_15 vdd gnd cell_6t
Xbit_r16_c242 bl_242 br_242 wl_16 vdd gnd cell_6t
Xbit_r17_c242 bl_242 br_242 wl_17 vdd gnd cell_6t
Xbit_r18_c242 bl_242 br_242 wl_18 vdd gnd cell_6t
Xbit_r19_c242 bl_242 br_242 wl_19 vdd gnd cell_6t
Xbit_r20_c242 bl_242 br_242 wl_20 vdd gnd cell_6t
Xbit_r21_c242 bl_242 br_242 wl_21 vdd gnd cell_6t
Xbit_r22_c242 bl_242 br_242 wl_22 vdd gnd cell_6t
Xbit_r23_c242 bl_242 br_242 wl_23 vdd gnd cell_6t
Xbit_r24_c242 bl_242 br_242 wl_24 vdd gnd cell_6t
Xbit_r25_c242 bl_242 br_242 wl_25 vdd gnd cell_6t
Xbit_r26_c242 bl_242 br_242 wl_26 vdd gnd cell_6t
Xbit_r27_c242 bl_242 br_242 wl_27 vdd gnd cell_6t
Xbit_r28_c242 bl_242 br_242 wl_28 vdd gnd cell_6t
Xbit_r29_c242 bl_242 br_242 wl_29 vdd gnd cell_6t
Xbit_r30_c242 bl_242 br_242 wl_30 vdd gnd cell_6t
Xbit_r31_c242 bl_242 br_242 wl_31 vdd gnd cell_6t
Xbit_r32_c242 bl_242 br_242 wl_32 vdd gnd cell_6t
Xbit_r33_c242 bl_242 br_242 wl_33 vdd gnd cell_6t
Xbit_r34_c242 bl_242 br_242 wl_34 vdd gnd cell_6t
Xbit_r35_c242 bl_242 br_242 wl_35 vdd gnd cell_6t
Xbit_r36_c242 bl_242 br_242 wl_36 vdd gnd cell_6t
Xbit_r37_c242 bl_242 br_242 wl_37 vdd gnd cell_6t
Xbit_r38_c242 bl_242 br_242 wl_38 vdd gnd cell_6t
Xbit_r39_c242 bl_242 br_242 wl_39 vdd gnd cell_6t
Xbit_r40_c242 bl_242 br_242 wl_40 vdd gnd cell_6t
Xbit_r41_c242 bl_242 br_242 wl_41 vdd gnd cell_6t
Xbit_r42_c242 bl_242 br_242 wl_42 vdd gnd cell_6t
Xbit_r43_c242 bl_242 br_242 wl_43 vdd gnd cell_6t
Xbit_r44_c242 bl_242 br_242 wl_44 vdd gnd cell_6t
Xbit_r45_c242 bl_242 br_242 wl_45 vdd gnd cell_6t
Xbit_r46_c242 bl_242 br_242 wl_46 vdd gnd cell_6t
Xbit_r47_c242 bl_242 br_242 wl_47 vdd gnd cell_6t
Xbit_r48_c242 bl_242 br_242 wl_48 vdd gnd cell_6t
Xbit_r49_c242 bl_242 br_242 wl_49 vdd gnd cell_6t
Xbit_r50_c242 bl_242 br_242 wl_50 vdd gnd cell_6t
Xbit_r51_c242 bl_242 br_242 wl_51 vdd gnd cell_6t
Xbit_r52_c242 bl_242 br_242 wl_52 vdd gnd cell_6t
Xbit_r53_c242 bl_242 br_242 wl_53 vdd gnd cell_6t
Xbit_r54_c242 bl_242 br_242 wl_54 vdd gnd cell_6t
Xbit_r55_c242 bl_242 br_242 wl_55 vdd gnd cell_6t
Xbit_r56_c242 bl_242 br_242 wl_56 vdd gnd cell_6t
Xbit_r57_c242 bl_242 br_242 wl_57 vdd gnd cell_6t
Xbit_r58_c242 bl_242 br_242 wl_58 vdd gnd cell_6t
Xbit_r59_c242 bl_242 br_242 wl_59 vdd gnd cell_6t
Xbit_r60_c242 bl_242 br_242 wl_60 vdd gnd cell_6t
Xbit_r61_c242 bl_242 br_242 wl_61 vdd gnd cell_6t
Xbit_r62_c242 bl_242 br_242 wl_62 vdd gnd cell_6t
Xbit_r63_c242 bl_242 br_242 wl_63 vdd gnd cell_6t
Xbit_r64_c242 bl_242 br_242 wl_64 vdd gnd cell_6t
Xbit_r65_c242 bl_242 br_242 wl_65 vdd gnd cell_6t
Xbit_r66_c242 bl_242 br_242 wl_66 vdd gnd cell_6t
Xbit_r67_c242 bl_242 br_242 wl_67 vdd gnd cell_6t
Xbit_r68_c242 bl_242 br_242 wl_68 vdd gnd cell_6t
Xbit_r69_c242 bl_242 br_242 wl_69 vdd gnd cell_6t
Xbit_r70_c242 bl_242 br_242 wl_70 vdd gnd cell_6t
Xbit_r71_c242 bl_242 br_242 wl_71 vdd gnd cell_6t
Xbit_r72_c242 bl_242 br_242 wl_72 vdd gnd cell_6t
Xbit_r73_c242 bl_242 br_242 wl_73 vdd gnd cell_6t
Xbit_r74_c242 bl_242 br_242 wl_74 vdd gnd cell_6t
Xbit_r75_c242 bl_242 br_242 wl_75 vdd gnd cell_6t
Xbit_r76_c242 bl_242 br_242 wl_76 vdd gnd cell_6t
Xbit_r77_c242 bl_242 br_242 wl_77 vdd gnd cell_6t
Xbit_r78_c242 bl_242 br_242 wl_78 vdd gnd cell_6t
Xbit_r79_c242 bl_242 br_242 wl_79 vdd gnd cell_6t
Xbit_r80_c242 bl_242 br_242 wl_80 vdd gnd cell_6t
Xbit_r81_c242 bl_242 br_242 wl_81 vdd gnd cell_6t
Xbit_r82_c242 bl_242 br_242 wl_82 vdd gnd cell_6t
Xbit_r83_c242 bl_242 br_242 wl_83 vdd gnd cell_6t
Xbit_r84_c242 bl_242 br_242 wl_84 vdd gnd cell_6t
Xbit_r85_c242 bl_242 br_242 wl_85 vdd gnd cell_6t
Xbit_r86_c242 bl_242 br_242 wl_86 vdd gnd cell_6t
Xbit_r87_c242 bl_242 br_242 wl_87 vdd gnd cell_6t
Xbit_r88_c242 bl_242 br_242 wl_88 vdd gnd cell_6t
Xbit_r89_c242 bl_242 br_242 wl_89 vdd gnd cell_6t
Xbit_r90_c242 bl_242 br_242 wl_90 vdd gnd cell_6t
Xbit_r91_c242 bl_242 br_242 wl_91 vdd gnd cell_6t
Xbit_r92_c242 bl_242 br_242 wl_92 vdd gnd cell_6t
Xbit_r93_c242 bl_242 br_242 wl_93 vdd gnd cell_6t
Xbit_r94_c242 bl_242 br_242 wl_94 vdd gnd cell_6t
Xbit_r95_c242 bl_242 br_242 wl_95 vdd gnd cell_6t
Xbit_r96_c242 bl_242 br_242 wl_96 vdd gnd cell_6t
Xbit_r97_c242 bl_242 br_242 wl_97 vdd gnd cell_6t
Xbit_r98_c242 bl_242 br_242 wl_98 vdd gnd cell_6t
Xbit_r99_c242 bl_242 br_242 wl_99 vdd gnd cell_6t
Xbit_r100_c242 bl_242 br_242 wl_100 vdd gnd cell_6t
Xbit_r101_c242 bl_242 br_242 wl_101 vdd gnd cell_6t
Xbit_r102_c242 bl_242 br_242 wl_102 vdd gnd cell_6t
Xbit_r103_c242 bl_242 br_242 wl_103 vdd gnd cell_6t
Xbit_r104_c242 bl_242 br_242 wl_104 vdd gnd cell_6t
Xbit_r105_c242 bl_242 br_242 wl_105 vdd gnd cell_6t
Xbit_r106_c242 bl_242 br_242 wl_106 vdd gnd cell_6t
Xbit_r107_c242 bl_242 br_242 wl_107 vdd gnd cell_6t
Xbit_r108_c242 bl_242 br_242 wl_108 vdd gnd cell_6t
Xbit_r109_c242 bl_242 br_242 wl_109 vdd gnd cell_6t
Xbit_r110_c242 bl_242 br_242 wl_110 vdd gnd cell_6t
Xbit_r111_c242 bl_242 br_242 wl_111 vdd gnd cell_6t
Xbit_r112_c242 bl_242 br_242 wl_112 vdd gnd cell_6t
Xbit_r113_c242 bl_242 br_242 wl_113 vdd gnd cell_6t
Xbit_r114_c242 bl_242 br_242 wl_114 vdd gnd cell_6t
Xbit_r115_c242 bl_242 br_242 wl_115 vdd gnd cell_6t
Xbit_r116_c242 bl_242 br_242 wl_116 vdd gnd cell_6t
Xbit_r117_c242 bl_242 br_242 wl_117 vdd gnd cell_6t
Xbit_r118_c242 bl_242 br_242 wl_118 vdd gnd cell_6t
Xbit_r119_c242 bl_242 br_242 wl_119 vdd gnd cell_6t
Xbit_r120_c242 bl_242 br_242 wl_120 vdd gnd cell_6t
Xbit_r121_c242 bl_242 br_242 wl_121 vdd gnd cell_6t
Xbit_r122_c242 bl_242 br_242 wl_122 vdd gnd cell_6t
Xbit_r123_c242 bl_242 br_242 wl_123 vdd gnd cell_6t
Xbit_r124_c242 bl_242 br_242 wl_124 vdd gnd cell_6t
Xbit_r125_c242 bl_242 br_242 wl_125 vdd gnd cell_6t
Xbit_r126_c242 bl_242 br_242 wl_126 vdd gnd cell_6t
Xbit_r127_c242 bl_242 br_242 wl_127 vdd gnd cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd cell_6t
Xbit_r1_c243 bl_243 br_243 wl_1 vdd gnd cell_6t
Xbit_r2_c243 bl_243 br_243 wl_2 vdd gnd cell_6t
Xbit_r3_c243 bl_243 br_243 wl_3 vdd gnd cell_6t
Xbit_r4_c243 bl_243 br_243 wl_4 vdd gnd cell_6t
Xbit_r5_c243 bl_243 br_243 wl_5 vdd gnd cell_6t
Xbit_r6_c243 bl_243 br_243 wl_6 vdd gnd cell_6t
Xbit_r7_c243 bl_243 br_243 wl_7 vdd gnd cell_6t
Xbit_r8_c243 bl_243 br_243 wl_8 vdd gnd cell_6t
Xbit_r9_c243 bl_243 br_243 wl_9 vdd gnd cell_6t
Xbit_r10_c243 bl_243 br_243 wl_10 vdd gnd cell_6t
Xbit_r11_c243 bl_243 br_243 wl_11 vdd gnd cell_6t
Xbit_r12_c243 bl_243 br_243 wl_12 vdd gnd cell_6t
Xbit_r13_c243 bl_243 br_243 wl_13 vdd gnd cell_6t
Xbit_r14_c243 bl_243 br_243 wl_14 vdd gnd cell_6t
Xbit_r15_c243 bl_243 br_243 wl_15 vdd gnd cell_6t
Xbit_r16_c243 bl_243 br_243 wl_16 vdd gnd cell_6t
Xbit_r17_c243 bl_243 br_243 wl_17 vdd gnd cell_6t
Xbit_r18_c243 bl_243 br_243 wl_18 vdd gnd cell_6t
Xbit_r19_c243 bl_243 br_243 wl_19 vdd gnd cell_6t
Xbit_r20_c243 bl_243 br_243 wl_20 vdd gnd cell_6t
Xbit_r21_c243 bl_243 br_243 wl_21 vdd gnd cell_6t
Xbit_r22_c243 bl_243 br_243 wl_22 vdd gnd cell_6t
Xbit_r23_c243 bl_243 br_243 wl_23 vdd gnd cell_6t
Xbit_r24_c243 bl_243 br_243 wl_24 vdd gnd cell_6t
Xbit_r25_c243 bl_243 br_243 wl_25 vdd gnd cell_6t
Xbit_r26_c243 bl_243 br_243 wl_26 vdd gnd cell_6t
Xbit_r27_c243 bl_243 br_243 wl_27 vdd gnd cell_6t
Xbit_r28_c243 bl_243 br_243 wl_28 vdd gnd cell_6t
Xbit_r29_c243 bl_243 br_243 wl_29 vdd gnd cell_6t
Xbit_r30_c243 bl_243 br_243 wl_30 vdd gnd cell_6t
Xbit_r31_c243 bl_243 br_243 wl_31 vdd gnd cell_6t
Xbit_r32_c243 bl_243 br_243 wl_32 vdd gnd cell_6t
Xbit_r33_c243 bl_243 br_243 wl_33 vdd gnd cell_6t
Xbit_r34_c243 bl_243 br_243 wl_34 vdd gnd cell_6t
Xbit_r35_c243 bl_243 br_243 wl_35 vdd gnd cell_6t
Xbit_r36_c243 bl_243 br_243 wl_36 vdd gnd cell_6t
Xbit_r37_c243 bl_243 br_243 wl_37 vdd gnd cell_6t
Xbit_r38_c243 bl_243 br_243 wl_38 vdd gnd cell_6t
Xbit_r39_c243 bl_243 br_243 wl_39 vdd gnd cell_6t
Xbit_r40_c243 bl_243 br_243 wl_40 vdd gnd cell_6t
Xbit_r41_c243 bl_243 br_243 wl_41 vdd gnd cell_6t
Xbit_r42_c243 bl_243 br_243 wl_42 vdd gnd cell_6t
Xbit_r43_c243 bl_243 br_243 wl_43 vdd gnd cell_6t
Xbit_r44_c243 bl_243 br_243 wl_44 vdd gnd cell_6t
Xbit_r45_c243 bl_243 br_243 wl_45 vdd gnd cell_6t
Xbit_r46_c243 bl_243 br_243 wl_46 vdd gnd cell_6t
Xbit_r47_c243 bl_243 br_243 wl_47 vdd gnd cell_6t
Xbit_r48_c243 bl_243 br_243 wl_48 vdd gnd cell_6t
Xbit_r49_c243 bl_243 br_243 wl_49 vdd gnd cell_6t
Xbit_r50_c243 bl_243 br_243 wl_50 vdd gnd cell_6t
Xbit_r51_c243 bl_243 br_243 wl_51 vdd gnd cell_6t
Xbit_r52_c243 bl_243 br_243 wl_52 vdd gnd cell_6t
Xbit_r53_c243 bl_243 br_243 wl_53 vdd gnd cell_6t
Xbit_r54_c243 bl_243 br_243 wl_54 vdd gnd cell_6t
Xbit_r55_c243 bl_243 br_243 wl_55 vdd gnd cell_6t
Xbit_r56_c243 bl_243 br_243 wl_56 vdd gnd cell_6t
Xbit_r57_c243 bl_243 br_243 wl_57 vdd gnd cell_6t
Xbit_r58_c243 bl_243 br_243 wl_58 vdd gnd cell_6t
Xbit_r59_c243 bl_243 br_243 wl_59 vdd gnd cell_6t
Xbit_r60_c243 bl_243 br_243 wl_60 vdd gnd cell_6t
Xbit_r61_c243 bl_243 br_243 wl_61 vdd gnd cell_6t
Xbit_r62_c243 bl_243 br_243 wl_62 vdd gnd cell_6t
Xbit_r63_c243 bl_243 br_243 wl_63 vdd gnd cell_6t
Xbit_r64_c243 bl_243 br_243 wl_64 vdd gnd cell_6t
Xbit_r65_c243 bl_243 br_243 wl_65 vdd gnd cell_6t
Xbit_r66_c243 bl_243 br_243 wl_66 vdd gnd cell_6t
Xbit_r67_c243 bl_243 br_243 wl_67 vdd gnd cell_6t
Xbit_r68_c243 bl_243 br_243 wl_68 vdd gnd cell_6t
Xbit_r69_c243 bl_243 br_243 wl_69 vdd gnd cell_6t
Xbit_r70_c243 bl_243 br_243 wl_70 vdd gnd cell_6t
Xbit_r71_c243 bl_243 br_243 wl_71 vdd gnd cell_6t
Xbit_r72_c243 bl_243 br_243 wl_72 vdd gnd cell_6t
Xbit_r73_c243 bl_243 br_243 wl_73 vdd gnd cell_6t
Xbit_r74_c243 bl_243 br_243 wl_74 vdd gnd cell_6t
Xbit_r75_c243 bl_243 br_243 wl_75 vdd gnd cell_6t
Xbit_r76_c243 bl_243 br_243 wl_76 vdd gnd cell_6t
Xbit_r77_c243 bl_243 br_243 wl_77 vdd gnd cell_6t
Xbit_r78_c243 bl_243 br_243 wl_78 vdd gnd cell_6t
Xbit_r79_c243 bl_243 br_243 wl_79 vdd gnd cell_6t
Xbit_r80_c243 bl_243 br_243 wl_80 vdd gnd cell_6t
Xbit_r81_c243 bl_243 br_243 wl_81 vdd gnd cell_6t
Xbit_r82_c243 bl_243 br_243 wl_82 vdd gnd cell_6t
Xbit_r83_c243 bl_243 br_243 wl_83 vdd gnd cell_6t
Xbit_r84_c243 bl_243 br_243 wl_84 vdd gnd cell_6t
Xbit_r85_c243 bl_243 br_243 wl_85 vdd gnd cell_6t
Xbit_r86_c243 bl_243 br_243 wl_86 vdd gnd cell_6t
Xbit_r87_c243 bl_243 br_243 wl_87 vdd gnd cell_6t
Xbit_r88_c243 bl_243 br_243 wl_88 vdd gnd cell_6t
Xbit_r89_c243 bl_243 br_243 wl_89 vdd gnd cell_6t
Xbit_r90_c243 bl_243 br_243 wl_90 vdd gnd cell_6t
Xbit_r91_c243 bl_243 br_243 wl_91 vdd gnd cell_6t
Xbit_r92_c243 bl_243 br_243 wl_92 vdd gnd cell_6t
Xbit_r93_c243 bl_243 br_243 wl_93 vdd gnd cell_6t
Xbit_r94_c243 bl_243 br_243 wl_94 vdd gnd cell_6t
Xbit_r95_c243 bl_243 br_243 wl_95 vdd gnd cell_6t
Xbit_r96_c243 bl_243 br_243 wl_96 vdd gnd cell_6t
Xbit_r97_c243 bl_243 br_243 wl_97 vdd gnd cell_6t
Xbit_r98_c243 bl_243 br_243 wl_98 vdd gnd cell_6t
Xbit_r99_c243 bl_243 br_243 wl_99 vdd gnd cell_6t
Xbit_r100_c243 bl_243 br_243 wl_100 vdd gnd cell_6t
Xbit_r101_c243 bl_243 br_243 wl_101 vdd gnd cell_6t
Xbit_r102_c243 bl_243 br_243 wl_102 vdd gnd cell_6t
Xbit_r103_c243 bl_243 br_243 wl_103 vdd gnd cell_6t
Xbit_r104_c243 bl_243 br_243 wl_104 vdd gnd cell_6t
Xbit_r105_c243 bl_243 br_243 wl_105 vdd gnd cell_6t
Xbit_r106_c243 bl_243 br_243 wl_106 vdd gnd cell_6t
Xbit_r107_c243 bl_243 br_243 wl_107 vdd gnd cell_6t
Xbit_r108_c243 bl_243 br_243 wl_108 vdd gnd cell_6t
Xbit_r109_c243 bl_243 br_243 wl_109 vdd gnd cell_6t
Xbit_r110_c243 bl_243 br_243 wl_110 vdd gnd cell_6t
Xbit_r111_c243 bl_243 br_243 wl_111 vdd gnd cell_6t
Xbit_r112_c243 bl_243 br_243 wl_112 vdd gnd cell_6t
Xbit_r113_c243 bl_243 br_243 wl_113 vdd gnd cell_6t
Xbit_r114_c243 bl_243 br_243 wl_114 vdd gnd cell_6t
Xbit_r115_c243 bl_243 br_243 wl_115 vdd gnd cell_6t
Xbit_r116_c243 bl_243 br_243 wl_116 vdd gnd cell_6t
Xbit_r117_c243 bl_243 br_243 wl_117 vdd gnd cell_6t
Xbit_r118_c243 bl_243 br_243 wl_118 vdd gnd cell_6t
Xbit_r119_c243 bl_243 br_243 wl_119 vdd gnd cell_6t
Xbit_r120_c243 bl_243 br_243 wl_120 vdd gnd cell_6t
Xbit_r121_c243 bl_243 br_243 wl_121 vdd gnd cell_6t
Xbit_r122_c243 bl_243 br_243 wl_122 vdd gnd cell_6t
Xbit_r123_c243 bl_243 br_243 wl_123 vdd gnd cell_6t
Xbit_r124_c243 bl_243 br_243 wl_124 vdd gnd cell_6t
Xbit_r125_c243 bl_243 br_243 wl_125 vdd gnd cell_6t
Xbit_r126_c243 bl_243 br_243 wl_126 vdd gnd cell_6t
Xbit_r127_c243 bl_243 br_243 wl_127 vdd gnd cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd cell_6t
Xbit_r1_c244 bl_244 br_244 wl_1 vdd gnd cell_6t
Xbit_r2_c244 bl_244 br_244 wl_2 vdd gnd cell_6t
Xbit_r3_c244 bl_244 br_244 wl_3 vdd gnd cell_6t
Xbit_r4_c244 bl_244 br_244 wl_4 vdd gnd cell_6t
Xbit_r5_c244 bl_244 br_244 wl_5 vdd gnd cell_6t
Xbit_r6_c244 bl_244 br_244 wl_6 vdd gnd cell_6t
Xbit_r7_c244 bl_244 br_244 wl_7 vdd gnd cell_6t
Xbit_r8_c244 bl_244 br_244 wl_8 vdd gnd cell_6t
Xbit_r9_c244 bl_244 br_244 wl_9 vdd gnd cell_6t
Xbit_r10_c244 bl_244 br_244 wl_10 vdd gnd cell_6t
Xbit_r11_c244 bl_244 br_244 wl_11 vdd gnd cell_6t
Xbit_r12_c244 bl_244 br_244 wl_12 vdd gnd cell_6t
Xbit_r13_c244 bl_244 br_244 wl_13 vdd gnd cell_6t
Xbit_r14_c244 bl_244 br_244 wl_14 vdd gnd cell_6t
Xbit_r15_c244 bl_244 br_244 wl_15 vdd gnd cell_6t
Xbit_r16_c244 bl_244 br_244 wl_16 vdd gnd cell_6t
Xbit_r17_c244 bl_244 br_244 wl_17 vdd gnd cell_6t
Xbit_r18_c244 bl_244 br_244 wl_18 vdd gnd cell_6t
Xbit_r19_c244 bl_244 br_244 wl_19 vdd gnd cell_6t
Xbit_r20_c244 bl_244 br_244 wl_20 vdd gnd cell_6t
Xbit_r21_c244 bl_244 br_244 wl_21 vdd gnd cell_6t
Xbit_r22_c244 bl_244 br_244 wl_22 vdd gnd cell_6t
Xbit_r23_c244 bl_244 br_244 wl_23 vdd gnd cell_6t
Xbit_r24_c244 bl_244 br_244 wl_24 vdd gnd cell_6t
Xbit_r25_c244 bl_244 br_244 wl_25 vdd gnd cell_6t
Xbit_r26_c244 bl_244 br_244 wl_26 vdd gnd cell_6t
Xbit_r27_c244 bl_244 br_244 wl_27 vdd gnd cell_6t
Xbit_r28_c244 bl_244 br_244 wl_28 vdd gnd cell_6t
Xbit_r29_c244 bl_244 br_244 wl_29 vdd gnd cell_6t
Xbit_r30_c244 bl_244 br_244 wl_30 vdd gnd cell_6t
Xbit_r31_c244 bl_244 br_244 wl_31 vdd gnd cell_6t
Xbit_r32_c244 bl_244 br_244 wl_32 vdd gnd cell_6t
Xbit_r33_c244 bl_244 br_244 wl_33 vdd gnd cell_6t
Xbit_r34_c244 bl_244 br_244 wl_34 vdd gnd cell_6t
Xbit_r35_c244 bl_244 br_244 wl_35 vdd gnd cell_6t
Xbit_r36_c244 bl_244 br_244 wl_36 vdd gnd cell_6t
Xbit_r37_c244 bl_244 br_244 wl_37 vdd gnd cell_6t
Xbit_r38_c244 bl_244 br_244 wl_38 vdd gnd cell_6t
Xbit_r39_c244 bl_244 br_244 wl_39 vdd gnd cell_6t
Xbit_r40_c244 bl_244 br_244 wl_40 vdd gnd cell_6t
Xbit_r41_c244 bl_244 br_244 wl_41 vdd gnd cell_6t
Xbit_r42_c244 bl_244 br_244 wl_42 vdd gnd cell_6t
Xbit_r43_c244 bl_244 br_244 wl_43 vdd gnd cell_6t
Xbit_r44_c244 bl_244 br_244 wl_44 vdd gnd cell_6t
Xbit_r45_c244 bl_244 br_244 wl_45 vdd gnd cell_6t
Xbit_r46_c244 bl_244 br_244 wl_46 vdd gnd cell_6t
Xbit_r47_c244 bl_244 br_244 wl_47 vdd gnd cell_6t
Xbit_r48_c244 bl_244 br_244 wl_48 vdd gnd cell_6t
Xbit_r49_c244 bl_244 br_244 wl_49 vdd gnd cell_6t
Xbit_r50_c244 bl_244 br_244 wl_50 vdd gnd cell_6t
Xbit_r51_c244 bl_244 br_244 wl_51 vdd gnd cell_6t
Xbit_r52_c244 bl_244 br_244 wl_52 vdd gnd cell_6t
Xbit_r53_c244 bl_244 br_244 wl_53 vdd gnd cell_6t
Xbit_r54_c244 bl_244 br_244 wl_54 vdd gnd cell_6t
Xbit_r55_c244 bl_244 br_244 wl_55 vdd gnd cell_6t
Xbit_r56_c244 bl_244 br_244 wl_56 vdd gnd cell_6t
Xbit_r57_c244 bl_244 br_244 wl_57 vdd gnd cell_6t
Xbit_r58_c244 bl_244 br_244 wl_58 vdd gnd cell_6t
Xbit_r59_c244 bl_244 br_244 wl_59 vdd gnd cell_6t
Xbit_r60_c244 bl_244 br_244 wl_60 vdd gnd cell_6t
Xbit_r61_c244 bl_244 br_244 wl_61 vdd gnd cell_6t
Xbit_r62_c244 bl_244 br_244 wl_62 vdd gnd cell_6t
Xbit_r63_c244 bl_244 br_244 wl_63 vdd gnd cell_6t
Xbit_r64_c244 bl_244 br_244 wl_64 vdd gnd cell_6t
Xbit_r65_c244 bl_244 br_244 wl_65 vdd gnd cell_6t
Xbit_r66_c244 bl_244 br_244 wl_66 vdd gnd cell_6t
Xbit_r67_c244 bl_244 br_244 wl_67 vdd gnd cell_6t
Xbit_r68_c244 bl_244 br_244 wl_68 vdd gnd cell_6t
Xbit_r69_c244 bl_244 br_244 wl_69 vdd gnd cell_6t
Xbit_r70_c244 bl_244 br_244 wl_70 vdd gnd cell_6t
Xbit_r71_c244 bl_244 br_244 wl_71 vdd gnd cell_6t
Xbit_r72_c244 bl_244 br_244 wl_72 vdd gnd cell_6t
Xbit_r73_c244 bl_244 br_244 wl_73 vdd gnd cell_6t
Xbit_r74_c244 bl_244 br_244 wl_74 vdd gnd cell_6t
Xbit_r75_c244 bl_244 br_244 wl_75 vdd gnd cell_6t
Xbit_r76_c244 bl_244 br_244 wl_76 vdd gnd cell_6t
Xbit_r77_c244 bl_244 br_244 wl_77 vdd gnd cell_6t
Xbit_r78_c244 bl_244 br_244 wl_78 vdd gnd cell_6t
Xbit_r79_c244 bl_244 br_244 wl_79 vdd gnd cell_6t
Xbit_r80_c244 bl_244 br_244 wl_80 vdd gnd cell_6t
Xbit_r81_c244 bl_244 br_244 wl_81 vdd gnd cell_6t
Xbit_r82_c244 bl_244 br_244 wl_82 vdd gnd cell_6t
Xbit_r83_c244 bl_244 br_244 wl_83 vdd gnd cell_6t
Xbit_r84_c244 bl_244 br_244 wl_84 vdd gnd cell_6t
Xbit_r85_c244 bl_244 br_244 wl_85 vdd gnd cell_6t
Xbit_r86_c244 bl_244 br_244 wl_86 vdd gnd cell_6t
Xbit_r87_c244 bl_244 br_244 wl_87 vdd gnd cell_6t
Xbit_r88_c244 bl_244 br_244 wl_88 vdd gnd cell_6t
Xbit_r89_c244 bl_244 br_244 wl_89 vdd gnd cell_6t
Xbit_r90_c244 bl_244 br_244 wl_90 vdd gnd cell_6t
Xbit_r91_c244 bl_244 br_244 wl_91 vdd gnd cell_6t
Xbit_r92_c244 bl_244 br_244 wl_92 vdd gnd cell_6t
Xbit_r93_c244 bl_244 br_244 wl_93 vdd gnd cell_6t
Xbit_r94_c244 bl_244 br_244 wl_94 vdd gnd cell_6t
Xbit_r95_c244 bl_244 br_244 wl_95 vdd gnd cell_6t
Xbit_r96_c244 bl_244 br_244 wl_96 vdd gnd cell_6t
Xbit_r97_c244 bl_244 br_244 wl_97 vdd gnd cell_6t
Xbit_r98_c244 bl_244 br_244 wl_98 vdd gnd cell_6t
Xbit_r99_c244 bl_244 br_244 wl_99 vdd gnd cell_6t
Xbit_r100_c244 bl_244 br_244 wl_100 vdd gnd cell_6t
Xbit_r101_c244 bl_244 br_244 wl_101 vdd gnd cell_6t
Xbit_r102_c244 bl_244 br_244 wl_102 vdd gnd cell_6t
Xbit_r103_c244 bl_244 br_244 wl_103 vdd gnd cell_6t
Xbit_r104_c244 bl_244 br_244 wl_104 vdd gnd cell_6t
Xbit_r105_c244 bl_244 br_244 wl_105 vdd gnd cell_6t
Xbit_r106_c244 bl_244 br_244 wl_106 vdd gnd cell_6t
Xbit_r107_c244 bl_244 br_244 wl_107 vdd gnd cell_6t
Xbit_r108_c244 bl_244 br_244 wl_108 vdd gnd cell_6t
Xbit_r109_c244 bl_244 br_244 wl_109 vdd gnd cell_6t
Xbit_r110_c244 bl_244 br_244 wl_110 vdd gnd cell_6t
Xbit_r111_c244 bl_244 br_244 wl_111 vdd gnd cell_6t
Xbit_r112_c244 bl_244 br_244 wl_112 vdd gnd cell_6t
Xbit_r113_c244 bl_244 br_244 wl_113 vdd gnd cell_6t
Xbit_r114_c244 bl_244 br_244 wl_114 vdd gnd cell_6t
Xbit_r115_c244 bl_244 br_244 wl_115 vdd gnd cell_6t
Xbit_r116_c244 bl_244 br_244 wl_116 vdd gnd cell_6t
Xbit_r117_c244 bl_244 br_244 wl_117 vdd gnd cell_6t
Xbit_r118_c244 bl_244 br_244 wl_118 vdd gnd cell_6t
Xbit_r119_c244 bl_244 br_244 wl_119 vdd gnd cell_6t
Xbit_r120_c244 bl_244 br_244 wl_120 vdd gnd cell_6t
Xbit_r121_c244 bl_244 br_244 wl_121 vdd gnd cell_6t
Xbit_r122_c244 bl_244 br_244 wl_122 vdd gnd cell_6t
Xbit_r123_c244 bl_244 br_244 wl_123 vdd gnd cell_6t
Xbit_r124_c244 bl_244 br_244 wl_124 vdd gnd cell_6t
Xbit_r125_c244 bl_244 br_244 wl_125 vdd gnd cell_6t
Xbit_r126_c244 bl_244 br_244 wl_126 vdd gnd cell_6t
Xbit_r127_c244 bl_244 br_244 wl_127 vdd gnd cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd cell_6t
Xbit_r1_c245 bl_245 br_245 wl_1 vdd gnd cell_6t
Xbit_r2_c245 bl_245 br_245 wl_2 vdd gnd cell_6t
Xbit_r3_c245 bl_245 br_245 wl_3 vdd gnd cell_6t
Xbit_r4_c245 bl_245 br_245 wl_4 vdd gnd cell_6t
Xbit_r5_c245 bl_245 br_245 wl_5 vdd gnd cell_6t
Xbit_r6_c245 bl_245 br_245 wl_6 vdd gnd cell_6t
Xbit_r7_c245 bl_245 br_245 wl_7 vdd gnd cell_6t
Xbit_r8_c245 bl_245 br_245 wl_8 vdd gnd cell_6t
Xbit_r9_c245 bl_245 br_245 wl_9 vdd gnd cell_6t
Xbit_r10_c245 bl_245 br_245 wl_10 vdd gnd cell_6t
Xbit_r11_c245 bl_245 br_245 wl_11 vdd gnd cell_6t
Xbit_r12_c245 bl_245 br_245 wl_12 vdd gnd cell_6t
Xbit_r13_c245 bl_245 br_245 wl_13 vdd gnd cell_6t
Xbit_r14_c245 bl_245 br_245 wl_14 vdd gnd cell_6t
Xbit_r15_c245 bl_245 br_245 wl_15 vdd gnd cell_6t
Xbit_r16_c245 bl_245 br_245 wl_16 vdd gnd cell_6t
Xbit_r17_c245 bl_245 br_245 wl_17 vdd gnd cell_6t
Xbit_r18_c245 bl_245 br_245 wl_18 vdd gnd cell_6t
Xbit_r19_c245 bl_245 br_245 wl_19 vdd gnd cell_6t
Xbit_r20_c245 bl_245 br_245 wl_20 vdd gnd cell_6t
Xbit_r21_c245 bl_245 br_245 wl_21 vdd gnd cell_6t
Xbit_r22_c245 bl_245 br_245 wl_22 vdd gnd cell_6t
Xbit_r23_c245 bl_245 br_245 wl_23 vdd gnd cell_6t
Xbit_r24_c245 bl_245 br_245 wl_24 vdd gnd cell_6t
Xbit_r25_c245 bl_245 br_245 wl_25 vdd gnd cell_6t
Xbit_r26_c245 bl_245 br_245 wl_26 vdd gnd cell_6t
Xbit_r27_c245 bl_245 br_245 wl_27 vdd gnd cell_6t
Xbit_r28_c245 bl_245 br_245 wl_28 vdd gnd cell_6t
Xbit_r29_c245 bl_245 br_245 wl_29 vdd gnd cell_6t
Xbit_r30_c245 bl_245 br_245 wl_30 vdd gnd cell_6t
Xbit_r31_c245 bl_245 br_245 wl_31 vdd gnd cell_6t
Xbit_r32_c245 bl_245 br_245 wl_32 vdd gnd cell_6t
Xbit_r33_c245 bl_245 br_245 wl_33 vdd gnd cell_6t
Xbit_r34_c245 bl_245 br_245 wl_34 vdd gnd cell_6t
Xbit_r35_c245 bl_245 br_245 wl_35 vdd gnd cell_6t
Xbit_r36_c245 bl_245 br_245 wl_36 vdd gnd cell_6t
Xbit_r37_c245 bl_245 br_245 wl_37 vdd gnd cell_6t
Xbit_r38_c245 bl_245 br_245 wl_38 vdd gnd cell_6t
Xbit_r39_c245 bl_245 br_245 wl_39 vdd gnd cell_6t
Xbit_r40_c245 bl_245 br_245 wl_40 vdd gnd cell_6t
Xbit_r41_c245 bl_245 br_245 wl_41 vdd gnd cell_6t
Xbit_r42_c245 bl_245 br_245 wl_42 vdd gnd cell_6t
Xbit_r43_c245 bl_245 br_245 wl_43 vdd gnd cell_6t
Xbit_r44_c245 bl_245 br_245 wl_44 vdd gnd cell_6t
Xbit_r45_c245 bl_245 br_245 wl_45 vdd gnd cell_6t
Xbit_r46_c245 bl_245 br_245 wl_46 vdd gnd cell_6t
Xbit_r47_c245 bl_245 br_245 wl_47 vdd gnd cell_6t
Xbit_r48_c245 bl_245 br_245 wl_48 vdd gnd cell_6t
Xbit_r49_c245 bl_245 br_245 wl_49 vdd gnd cell_6t
Xbit_r50_c245 bl_245 br_245 wl_50 vdd gnd cell_6t
Xbit_r51_c245 bl_245 br_245 wl_51 vdd gnd cell_6t
Xbit_r52_c245 bl_245 br_245 wl_52 vdd gnd cell_6t
Xbit_r53_c245 bl_245 br_245 wl_53 vdd gnd cell_6t
Xbit_r54_c245 bl_245 br_245 wl_54 vdd gnd cell_6t
Xbit_r55_c245 bl_245 br_245 wl_55 vdd gnd cell_6t
Xbit_r56_c245 bl_245 br_245 wl_56 vdd gnd cell_6t
Xbit_r57_c245 bl_245 br_245 wl_57 vdd gnd cell_6t
Xbit_r58_c245 bl_245 br_245 wl_58 vdd gnd cell_6t
Xbit_r59_c245 bl_245 br_245 wl_59 vdd gnd cell_6t
Xbit_r60_c245 bl_245 br_245 wl_60 vdd gnd cell_6t
Xbit_r61_c245 bl_245 br_245 wl_61 vdd gnd cell_6t
Xbit_r62_c245 bl_245 br_245 wl_62 vdd gnd cell_6t
Xbit_r63_c245 bl_245 br_245 wl_63 vdd gnd cell_6t
Xbit_r64_c245 bl_245 br_245 wl_64 vdd gnd cell_6t
Xbit_r65_c245 bl_245 br_245 wl_65 vdd gnd cell_6t
Xbit_r66_c245 bl_245 br_245 wl_66 vdd gnd cell_6t
Xbit_r67_c245 bl_245 br_245 wl_67 vdd gnd cell_6t
Xbit_r68_c245 bl_245 br_245 wl_68 vdd gnd cell_6t
Xbit_r69_c245 bl_245 br_245 wl_69 vdd gnd cell_6t
Xbit_r70_c245 bl_245 br_245 wl_70 vdd gnd cell_6t
Xbit_r71_c245 bl_245 br_245 wl_71 vdd gnd cell_6t
Xbit_r72_c245 bl_245 br_245 wl_72 vdd gnd cell_6t
Xbit_r73_c245 bl_245 br_245 wl_73 vdd gnd cell_6t
Xbit_r74_c245 bl_245 br_245 wl_74 vdd gnd cell_6t
Xbit_r75_c245 bl_245 br_245 wl_75 vdd gnd cell_6t
Xbit_r76_c245 bl_245 br_245 wl_76 vdd gnd cell_6t
Xbit_r77_c245 bl_245 br_245 wl_77 vdd gnd cell_6t
Xbit_r78_c245 bl_245 br_245 wl_78 vdd gnd cell_6t
Xbit_r79_c245 bl_245 br_245 wl_79 vdd gnd cell_6t
Xbit_r80_c245 bl_245 br_245 wl_80 vdd gnd cell_6t
Xbit_r81_c245 bl_245 br_245 wl_81 vdd gnd cell_6t
Xbit_r82_c245 bl_245 br_245 wl_82 vdd gnd cell_6t
Xbit_r83_c245 bl_245 br_245 wl_83 vdd gnd cell_6t
Xbit_r84_c245 bl_245 br_245 wl_84 vdd gnd cell_6t
Xbit_r85_c245 bl_245 br_245 wl_85 vdd gnd cell_6t
Xbit_r86_c245 bl_245 br_245 wl_86 vdd gnd cell_6t
Xbit_r87_c245 bl_245 br_245 wl_87 vdd gnd cell_6t
Xbit_r88_c245 bl_245 br_245 wl_88 vdd gnd cell_6t
Xbit_r89_c245 bl_245 br_245 wl_89 vdd gnd cell_6t
Xbit_r90_c245 bl_245 br_245 wl_90 vdd gnd cell_6t
Xbit_r91_c245 bl_245 br_245 wl_91 vdd gnd cell_6t
Xbit_r92_c245 bl_245 br_245 wl_92 vdd gnd cell_6t
Xbit_r93_c245 bl_245 br_245 wl_93 vdd gnd cell_6t
Xbit_r94_c245 bl_245 br_245 wl_94 vdd gnd cell_6t
Xbit_r95_c245 bl_245 br_245 wl_95 vdd gnd cell_6t
Xbit_r96_c245 bl_245 br_245 wl_96 vdd gnd cell_6t
Xbit_r97_c245 bl_245 br_245 wl_97 vdd gnd cell_6t
Xbit_r98_c245 bl_245 br_245 wl_98 vdd gnd cell_6t
Xbit_r99_c245 bl_245 br_245 wl_99 vdd gnd cell_6t
Xbit_r100_c245 bl_245 br_245 wl_100 vdd gnd cell_6t
Xbit_r101_c245 bl_245 br_245 wl_101 vdd gnd cell_6t
Xbit_r102_c245 bl_245 br_245 wl_102 vdd gnd cell_6t
Xbit_r103_c245 bl_245 br_245 wl_103 vdd gnd cell_6t
Xbit_r104_c245 bl_245 br_245 wl_104 vdd gnd cell_6t
Xbit_r105_c245 bl_245 br_245 wl_105 vdd gnd cell_6t
Xbit_r106_c245 bl_245 br_245 wl_106 vdd gnd cell_6t
Xbit_r107_c245 bl_245 br_245 wl_107 vdd gnd cell_6t
Xbit_r108_c245 bl_245 br_245 wl_108 vdd gnd cell_6t
Xbit_r109_c245 bl_245 br_245 wl_109 vdd gnd cell_6t
Xbit_r110_c245 bl_245 br_245 wl_110 vdd gnd cell_6t
Xbit_r111_c245 bl_245 br_245 wl_111 vdd gnd cell_6t
Xbit_r112_c245 bl_245 br_245 wl_112 vdd gnd cell_6t
Xbit_r113_c245 bl_245 br_245 wl_113 vdd gnd cell_6t
Xbit_r114_c245 bl_245 br_245 wl_114 vdd gnd cell_6t
Xbit_r115_c245 bl_245 br_245 wl_115 vdd gnd cell_6t
Xbit_r116_c245 bl_245 br_245 wl_116 vdd gnd cell_6t
Xbit_r117_c245 bl_245 br_245 wl_117 vdd gnd cell_6t
Xbit_r118_c245 bl_245 br_245 wl_118 vdd gnd cell_6t
Xbit_r119_c245 bl_245 br_245 wl_119 vdd gnd cell_6t
Xbit_r120_c245 bl_245 br_245 wl_120 vdd gnd cell_6t
Xbit_r121_c245 bl_245 br_245 wl_121 vdd gnd cell_6t
Xbit_r122_c245 bl_245 br_245 wl_122 vdd gnd cell_6t
Xbit_r123_c245 bl_245 br_245 wl_123 vdd gnd cell_6t
Xbit_r124_c245 bl_245 br_245 wl_124 vdd gnd cell_6t
Xbit_r125_c245 bl_245 br_245 wl_125 vdd gnd cell_6t
Xbit_r126_c245 bl_245 br_245 wl_126 vdd gnd cell_6t
Xbit_r127_c245 bl_245 br_245 wl_127 vdd gnd cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd cell_6t
Xbit_r1_c246 bl_246 br_246 wl_1 vdd gnd cell_6t
Xbit_r2_c246 bl_246 br_246 wl_2 vdd gnd cell_6t
Xbit_r3_c246 bl_246 br_246 wl_3 vdd gnd cell_6t
Xbit_r4_c246 bl_246 br_246 wl_4 vdd gnd cell_6t
Xbit_r5_c246 bl_246 br_246 wl_5 vdd gnd cell_6t
Xbit_r6_c246 bl_246 br_246 wl_6 vdd gnd cell_6t
Xbit_r7_c246 bl_246 br_246 wl_7 vdd gnd cell_6t
Xbit_r8_c246 bl_246 br_246 wl_8 vdd gnd cell_6t
Xbit_r9_c246 bl_246 br_246 wl_9 vdd gnd cell_6t
Xbit_r10_c246 bl_246 br_246 wl_10 vdd gnd cell_6t
Xbit_r11_c246 bl_246 br_246 wl_11 vdd gnd cell_6t
Xbit_r12_c246 bl_246 br_246 wl_12 vdd gnd cell_6t
Xbit_r13_c246 bl_246 br_246 wl_13 vdd gnd cell_6t
Xbit_r14_c246 bl_246 br_246 wl_14 vdd gnd cell_6t
Xbit_r15_c246 bl_246 br_246 wl_15 vdd gnd cell_6t
Xbit_r16_c246 bl_246 br_246 wl_16 vdd gnd cell_6t
Xbit_r17_c246 bl_246 br_246 wl_17 vdd gnd cell_6t
Xbit_r18_c246 bl_246 br_246 wl_18 vdd gnd cell_6t
Xbit_r19_c246 bl_246 br_246 wl_19 vdd gnd cell_6t
Xbit_r20_c246 bl_246 br_246 wl_20 vdd gnd cell_6t
Xbit_r21_c246 bl_246 br_246 wl_21 vdd gnd cell_6t
Xbit_r22_c246 bl_246 br_246 wl_22 vdd gnd cell_6t
Xbit_r23_c246 bl_246 br_246 wl_23 vdd gnd cell_6t
Xbit_r24_c246 bl_246 br_246 wl_24 vdd gnd cell_6t
Xbit_r25_c246 bl_246 br_246 wl_25 vdd gnd cell_6t
Xbit_r26_c246 bl_246 br_246 wl_26 vdd gnd cell_6t
Xbit_r27_c246 bl_246 br_246 wl_27 vdd gnd cell_6t
Xbit_r28_c246 bl_246 br_246 wl_28 vdd gnd cell_6t
Xbit_r29_c246 bl_246 br_246 wl_29 vdd gnd cell_6t
Xbit_r30_c246 bl_246 br_246 wl_30 vdd gnd cell_6t
Xbit_r31_c246 bl_246 br_246 wl_31 vdd gnd cell_6t
Xbit_r32_c246 bl_246 br_246 wl_32 vdd gnd cell_6t
Xbit_r33_c246 bl_246 br_246 wl_33 vdd gnd cell_6t
Xbit_r34_c246 bl_246 br_246 wl_34 vdd gnd cell_6t
Xbit_r35_c246 bl_246 br_246 wl_35 vdd gnd cell_6t
Xbit_r36_c246 bl_246 br_246 wl_36 vdd gnd cell_6t
Xbit_r37_c246 bl_246 br_246 wl_37 vdd gnd cell_6t
Xbit_r38_c246 bl_246 br_246 wl_38 vdd gnd cell_6t
Xbit_r39_c246 bl_246 br_246 wl_39 vdd gnd cell_6t
Xbit_r40_c246 bl_246 br_246 wl_40 vdd gnd cell_6t
Xbit_r41_c246 bl_246 br_246 wl_41 vdd gnd cell_6t
Xbit_r42_c246 bl_246 br_246 wl_42 vdd gnd cell_6t
Xbit_r43_c246 bl_246 br_246 wl_43 vdd gnd cell_6t
Xbit_r44_c246 bl_246 br_246 wl_44 vdd gnd cell_6t
Xbit_r45_c246 bl_246 br_246 wl_45 vdd gnd cell_6t
Xbit_r46_c246 bl_246 br_246 wl_46 vdd gnd cell_6t
Xbit_r47_c246 bl_246 br_246 wl_47 vdd gnd cell_6t
Xbit_r48_c246 bl_246 br_246 wl_48 vdd gnd cell_6t
Xbit_r49_c246 bl_246 br_246 wl_49 vdd gnd cell_6t
Xbit_r50_c246 bl_246 br_246 wl_50 vdd gnd cell_6t
Xbit_r51_c246 bl_246 br_246 wl_51 vdd gnd cell_6t
Xbit_r52_c246 bl_246 br_246 wl_52 vdd gnd cell_6t
Xbit_r53_c246 bl_246 br_246 wl_53 vdd gnd cell_6t
Xbit_r54_c246 bl_246 br_246 wl_54 vdd gnd cell_6t
Xbit_r55_c246 bl_246 br_246 wl_55 vdd gnd cell_6t
Xbit_r56_c246 bl_246 br_246 wl_56 vdd gnd cell_6t
Xbit_r57_c246 bl_246 br_246 wl_57 vdd gnd cell_6t
Xbit_r58_c246 bl_246 br_246 wl_58 vdd gnd cell_6t
Xbit_r59_c246 bl_246 br_246 wl_59 vdd gnd cell_6t
Xbit_r60_c246 bl_246 br_246 wl_60 vdd gnd cell_6t
Xbit_r61_c246 bl_246 br_246 wl_61 vdd gnd cell_6t
Xbit_r62_c246 bl_246 br_246 wl_62 vdd gnd cell_6t
Xbit_r63_c246 bl_246 br_246 wl_63 vdd gnd cell_6t
Xbit_r64_c246 bl_246 br_246 wl_64 vdd gnd cell_6t
Xbit_r65_c246 bl_246 br_246 wl_65 vdd gnd cell_6t
Xbit_r66_c246 bl_246 br_246 wl_66 vdd gnd cell_6t
Xbit_r67_c246 bl_246 br_246 wl_67 vdd gnd cell_6t
Xbit_r68_c246 bl_246 br_246 wl_68 vdd gnd cell_6t
Xbit_r69_c246 bl_246 br_246 wl_69 vdd gnd cell_6t
Xbit_r70_c246 bl_246 br_246 wl_70 vdd gnd cell_6t
Xbit_r71_c246 bl_246 br_246 wl_71 vdd gnd cell_6t
Xbit_r72_c246 bl_246 br_246 wl_72 vdd gnd cell_6t
Xbit_r73_c246 bl_246 br_246 wl_73 vdd gnd cell_6t
Xbit_r74_c246 bl_246 br_246 wl_74 vdd gnd cell_6t
Xbit_r75_c246 bl_246 br_246 wl_75 vdd gnd cell_6t
Xbit_r76_c246 bl_246 br_246 wl_76 vdd gnd cell_6t
Xbit_r77_c246 bl_246 br_246 wl_77 vdd gnd cell_6t
Xbit_r78_c246 bl_246 br_246 wl_78 vdd gnd cell_6t
Xbit_r79_c246 bl_246 br_246 wl_79 vdd gnd cell_6t
Xbit_r80_c246 bl_246 br_246 wl_80 vdd gnd cell_6t
Xbit_r81_c246 bl_246 br_246 wl_81 vdd gnd cell_6t
Xbit_r82_c246 bl_246 br_246 wl_82 vdd gnd cell_6t
Xbit_r83_c246 bl_246 br_246 wl_83 vdd gnd cell_6t
Xbit_r84_c246 bl_246 br_246 wl_84 vdd gnd cell_6t
Xbit_r85_c246 bl_246 br_246 wl_85 vdd gnd cell_6t
Xbit_r86_c246 bl_246 br_246 wl_86 vdd gnd cell_6t
Xbit_r87_c246 bl_246 br_246 wl_87 vdd gnd cell_6t
Xbit_r88_c246 bl_246 br_246 wl_88 vdd gnd cell_6t
Xbit_r89_c246 bl_246 br_246 wl_89 vdd gnd cell_6t
Xbit_r90_c246 bl_246 br_246 wl_90 vdd gnd cell_6t
Xbit_r91_c246 bl_246 br_246 wl_91 vdd gnd cell_6t
Xbit_r92_c246 bl_246 br_246 wl_92 vdd gnd cell_6t
Xbit_r93_c246 bl_246 br_246 wl_93 vdd gnd cell_6t
Xbit_r94_c246 bl_246 br_246 wl_94 vdd gnd cell_6t
Xbit_r95_c246 bl_246 br_246 wl_95 vdd gnd cell_6t
Xbit_r96_c246 bl_246 br_246 wl_96 vdd gnd cell_6t
Xbit_r97_c246 bl_246 br_246 wl_97 vdd gnd cell_6t
Xbit_r98_c246 bl_246 br_246 wl_98 vdd gnd cell_6t
Xbit_r99_c246 bl_246 br_246 wl_99 vdd gnd cell_6t
Xbit_r100_c246 bl_246 br_246 wl_100 vdd gnd cell_6t
Xbit_r101_c246 bl_246 br_246 wl_101 vdd gnd cell_6t
Xbit_r102_c246 bl_246 br_246 wl_102 vdd gnd cell_6t
Xbit_r103_c246 bl_246 br_246 wl_103 vdd gnd cell_6t
Xbit_r104_c246 bl_246 br_246 wl_104 vdd gnd cell_6t
Xbit_r105_c246 bl_246 br_246 wl_105 vdd gnd cell_6t
Xbit_r106_c246 bl_246 br_246 wl_106 vdd gnd cell_6t
Xbit_r107_c246 bl_246 br_246 wl_107 vdd gnd cell_6t
Xbit_r108_c246 bl_246 br_246 wl_108 vdd gnd cell_6t
Xbit_r109_c246 bl_246 br_246 wl_109 vdd gnd cell_6t
Xbit_r110_c246 bl_246 br_246 wl_110 vdd gnd cell_6t
Xbit_r111_c246 bl_246 br_246 wl_111 vdd gnd cell_6t
Xbit_r112_c246 bl_246 br_246 wl_112 vdd gnd cell_6t
Xbit_r113_c246 bl_246 br_246 wl_113 vdd gnd cell_6t
Xbit_r114_c246 bl_246 br_246 wl_114 vdd gnd cell_6t
Xbit_r115_c246 bl_246 br_246 wl_115 vdd gnd cell_6t
Xbit_r116_c246 bl_246 br_246 wl_116 vdd gnd cell_6t
Xbit_r117_c246 bl_246 br_246 wl_117 vdd gnd cell_6t
Xbit_r118_c246 bl_246 br_246 wl_118 vdd gnd cell_6t
Xbit_r119_c246 bl_246 br_246 wl_119 vdd gnd cell_6t
Xbit_r120_c246 bl_246 br_246 wl_120 vdd gnd cell_6t
Xbit_r121_c246 bl_246 br_246 wl_121 vdd gnd cell_6t
Xbit_r122_c246 bl_246 br_246 wl_122 vdd gnd cell_6t
Xbit_r123_c246 bl_246 br_246 wl_123 vdd gnd cell_6t
Xbit_r124_c246 bl_246 br_246 wl_124 vdd gnd cell_6t
Xbit_r125_c246 bl_246 br_246 wl_125 vdd gnd cell_6t
Xbit_r126_c246 bl_246 br_246 wl_126 vdd gnd cell_6t
Xbit_r127_c246 bl_246 br_246 wl_127 vdd gnd cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd cell_6t
Xbit_r1_c247 bl_247 br_247 wl_1 vdd gnd cell_6t
Xbit_r2_c247 bl_247 br_247 wl_2 vdd gnd cell_6t
Xbit_r3_c247 bl_247 br_247 wl_3 vdd gnd cell_6t
Xbit_r4_c247 bl_247 br_247 wl_4 vdd gnd cell_6t
Xbit_r5_c247 bl_247 br_247 wl_5 vdd gnd cell_6t
Xbit_r6_c247 bl_247 br_247 wl_6 vdd gnd cell_6t
Xbit_r7_c247 bl_247 br_247 wl_7 vdd gnd cell_6t
Xbit_r8_c247 bl_247 br_247 wl_8 vdd gnd cell_6t
Xbit_r9_c247 bl_247 br_247 wl_9 vdd gnd cell_6t
Xbit_r10_c247 bl_247 br_247 wl_10 vdd gnd cell_6t
Xbit_r11_c247 bl_247 br_247 wl_11 vdd gnd cell_6t
Xbit_r12_c247 bl_247 br_247 wl_12 vdd gnd cell_6t
Xbit_r13_c247 bl_247 br_247 wl_13 vdd gnd cell_6t
Xbit_r14_c247 bl_247 br_247 wl_14 vdd gnd cell_6t
Xbit_r15_c247 bl_247 br_247 wl_15 vdd gnd cell_6t
Xbit_r16_c247 bl_247 br_247 wl_16 vdd gnd cell_6t
Xbit_r17_c247 bl_247 br_247 wl_17 vdd gnd cell_6t
Xbit_r18_c247 bl_247 br_247 wl_18 vdd gnd cell_6t
Xbit_r19_c247 bl_247 br_247 wl_19 vdd gnd cell_6t
Xbit_r20_c247 bl_247 br_247 wl_20 vdd gnd cell_6t
Xbit_r21_c247 bl_247 br_247 wl_21 vdd gnd cell_6t
Xbit_r22_c247 bl_247 br_247 wl_22 vdd gnd cell_6t
Xbit_r23_c247 bl_247 br_247 wl_23 vdd gnd cell_6t
Xbit_r24_c247 bl_247 br_247 wl_24 vdd gnd cell_6t
Xbit_r25_c247 bl_247 br_247 wl_25 vdd gnd cell_6t
Xbit_r26_c247 bl_247 br_247 wl_26 vdd gnd cell_6t
Xbit_r27_c247 bl_247 br_247 wl_27 vdd gnd cell_6t
Xbit_r28_c247 bl_247 br_247 wl_28 vdd gnd cell_6t
Xbit_r29_c247 bl_247 br_247 wl_29 vdd gnd cell_6t
Xbit_r30_c247 bl_247 br_247 wl_30 vdd gnd cell_6t
Xbit_r31_c247 bl_247 br_247 wl_31 vdd gnd cell_6t
Xbit_r32_c247 bl_247 br_247 wl_32 vdd gnd cell_6t
Xbit_r33_c247 bl_247 br_247 wl_33 vdd gnd cell_6t
Xbit_r34_c247 bl_247 br_247 wl_34 vdd gnd cell_6t
Xbit_r35_c247 bl_247 br_247 wl_35 vdd gnd cell_6t
Xbit_r36_c247 bl_247 br_247 wl_36 vdd gnd cell_6t
Xbit_r37_c247 bl_247 br_247 wl_37 vdd gnd cell_6t
Xbit_r38_c247 bl_247 br_247 wl_38 vdd gnd cell_6t
Xbit_r39_c247 bl_247 br_247 wl_39 vdd gnd cell_6t
Xbit_r40_c247 bl_247 br_247 wl_40 vdd gnd cell_6t
Xbit_r41_c247 bl_247 br_247 wl_41 vdd gnd cell_6t
Xbit_r42_c247 bl_247 br_247 wl_42 vdd gnd cell_6t
Xbit_r43_c247 bl_247 br_247 wl_43 vdd gnd cell_6t
Xbit_r44_c247 bl_247 br_247 wl_44 vdd gnd cell_6t
Xbit_r45_c247 bl_247 br_247 wl_45 vdd gnd cell_6t
Xbit_r46_c247 bl_247 br_247 wl_46 vdd gnd cell_6t
Xbit_r47_c247 bl_247 br_247 wl_47 vdd gnd cell_6t
Xbit_r48_c247 bl_247 br_247 wl_48 vdd gnd cell_6t
Xbit_r49_c247 bl_247 br_247 wl_49 vdd gnd cell_6t
Xbit_r50_c247 bl_247 br_247 wl_50 vdd gnd cell_6t
Xbit_r51_c247 bl_247 br_247 wl_51 vdd gnd cell_6t
Xbit_r52_c247 bl_247 br_247 wl_52 vdd gnd cell_6t
Xbit_r53_c247 bl_247 br_247 wl_53 vdd gnd cell_6t
Xbit_r54_c247 bl_247 br_247 wl_54 vdd gnd cell_6t
Xbit_r55_c247 bl_247 br_247 wl_55 vdd gnd cell_6t
Xbit_r56_c247 bl_247 br_247 wl_56 vdd gnd cell_6t
Xbit_r57_c247 bl_247 br_247 wl_57 vdd gnd cell_6t
Xbit_r58_c247 bl_247 br_247 wl_58 vdd gnd cell_6t
Xbit_r59_c247 bl_247 br_247 wl_59 vdd gnd cell_6t
Xbit_r60_c247 bl_247 br_247 wl_60 vdd gnd cell_6t
Xbit_r61_c247 bl_247 br_247 wl_61 vdd gnd cell_6t
Xbit_r62_c247 bl_247 br_247 wl_62 vdd gnd cell_6t
Xbit_r63_c247 bl_247 br_247 wl_63 vdd gnd cell_6t
Xbit_r64_c247 bl_247 br_247 wl_64 vdd gnd cell_6t
Xbit_r65_c247 bl_247 br_247 wl_65 vdd gnd cell_6t
Xbit_r66_c247 bl_247 br_247 wl_66 vdd gnd cell_6t
Xbit_r67_c247 bl_247 br_247 wl_67 vdd gnd cell_6t
Xbit_r68_c247 bl_247 br_247 wl_68 vdd gnd cell_6t
Xbit_r69_c247 bl_247 br_247 wl_69 vdd gnd cell_6t
Xbit_r70_c247 bl_247 br_247 wl_70 vdd gnd cell_6t
Xbit_r71_c247 bl_247 br_247 wl_71 vdd gnd cell_6t
Xbit_r72_c247 bl_247 br_247 wl_72 vdd gnd cell_6t
Xbit_r73_c247 bl_247 br_247 wl_73 vdd gnd cell_6t
Xbit_r74_c247 bl_247 br_247 wl_74 vdd gnd cell_6t
Xbit_r75_c247 bl_247 br_247 wl_75 vdd gnd cell_6t
Xbit_r76_c247 bl_247 br_247 wl_76 vdd gnd cell_6t
Xbit_r77_c247 bl_247 br_247 wl_77 vdd gnd cell_6t
Xbit_r78_c247 bl_247 br_247 wl_78 vdd gnd cell_6t
Xbit_r79_c247 bl_247 br_247 wl_79 vdd gnd cell_6t
Xbit_r80_c247 bl_247 br_247 wl_80 vdd gnd cell_6t
Xbit_r81_c247 bl_247 br_247 wl_81 vdd gnd cell_6t
Xbit_r82_c247 bl_247 br_247 wl_82 vdd gnd cell_6t
Xbit_r83_c247 bl_247 br_247 wl_83 vdd gnd cell_6t
Xbit_r84_c247 bl_247 br_247 wl_84 vdd gnd cell_6t
Xbit_r85_c247 bl_247 br_247 wl_85 vdd gnd cell_6t
Xbit_r86_c247 bl_247 br_247 wl_86 vdd gnd cell_6t
Xbit_r87_c247 bl_247 br_247 wl_87 vdd gnd cell_6t
Xbit_r88_c247 bl_247 br_247 wl_88 vdd gnd cell_6t
Xbit_r89_c247 bl_247 br_247 wl_89 vdd gnd cell_6t
Xbit_r90_c247 bl_247 br_247 wl_90 vdd gnd cell_6t
Xbit_r91_c247 bl_247 br_247 wl_91 vdd gnd cell_6t
Xbit_r92_c247 bl_247 br_247 wl_92 vdd gnd cell_6t
Xbit_r93_c247 bl_247 br_247 wl_93 vdd gnd cell_6t
Xbit_r94_c247 bl_247 br_247 wl_94 vdd gnd cell_6t
Xbit_r95_c247 bl_247 br_247 wl_95 vdd gnd cell_6t
Xbit_r96_c247 bl_247 br_247 wl_96 vdd gnd cell_6t
Xbit_r97_c247 bl_247 br_247 wl_97 vdd gnd cell_6t
Xbit_r98_c247 bl_247 br_247 wl_98 vdd gnd cell_6t
Xbit_r99_c247 bl_247 br_247 wl_99 vdd gnd cell_6t
Xbit_r100_c247 bl_247 br_247 wl_100 vdd gnd cell_6t
Xbit_r101_c247 bl_247 br_247 wl_101 vdd gnd cell_6t
Xbit_r102_c247 bl_247 br_247 wl_102 vdd gnd cell_6t
Xbit_r103_c247 bl_247 br_247 wl_103 vdd gnd cell_6t
Xbit_r104_c247 bl_247 br_247 wl_104 vdd gnd cell_6t
Xbit_r105_c247 bl_247 br_247 wl_105 vdd gnd cell_6t
Xbit_r106_c247 bl_247 br_247 wl_106 vdd gnd cell_6t
Xbit_r107_c247 bl_247 br_247 wl_107 vdd gnd cell_6t
Xbit_r108_c247 bl_247 br_247 wl_108 vdd gnd cell_6t
Xbit_r109_c247 bl_247 br_247 wl_109 vdd gnd cell_6t
Xbit_r110_c247 bl_247 br_247 wl_110 vdd gnd cell_6t
Xbit_r111_c247 bl_247 br_247 wl_111 vdd gnd cell_6t
Xbit_r112_c247 bl_247 br_247 wl_112 vdd gnd cell_6t
Xbit_r113_c247 bl_247 br_247 wl_113 vdd gnd cell_6t
Xbit_r114_c247 bl_247 br_247 wl_114 vdd gnd cell_6t
Xbit_r115_c247 bl_247 br_247 wl_115 vdd gnd cell_6t
Xbit_r116_c247 bl_247 br_247 wl_116 vdd gnd cell_6t
Xbit_r117_c247 bl_247 br_247 wl_117 vdd gnd cell_6t
Xbit_r118_c247 bl_247 br_247 wl_118 vdd gnd cell_6t
Xbit_r119_c247 bl_247 br_247 wl_119 vdd gnd cell_6t
Xbit_r120_c247 bl_247 br_247 wl_120 vdd gnd cell_6t
Xbit_r121_c247 bl_247 br_247 wl_121 vdd gnd cell_6t
Xbit_r122_c247 bl_247 br_247 wl_122 vdd gnd cell_6t
Xbit_r123_c247 bl_247 br_247 wl_123 vdd gnd cell_6t
Xbit_r124_c247 bl_247 br_247 wl_124 vdd gnd cell_6t
Xbit_r125_c247 bl_247 br_247 wl_125 vdd gnd cell_6t
Xbit_r126_c247 bl_247 br_247 wl_126 vdd gnd cell_6t
Xbit_r127_c247 bl_247 br_247 wl_127 vdd gnd cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd cell_6t
Xbit_r1_c248 bl_248 br_248 wl_1 vdd gnd cell_6t
Xbit_r2_c248 bl_248 br_248 wl_2 vdd gnd cell_6t
Xbit_r3_c248 bl_248 br_248 wl_3 vdd gnd cell_6t
Xbit_r4_c248 bl_248 br_248 wl_4 vdd gnd cell_6t
Xbit_r5_c248 bl_248 br_248 wl_5 vdd gnd cell_6t
Xbit_r6_c248 bl_248 br_248 wl_6 vdd gnd cell_6t
Xbit_r7_c248 bl_248 br_248 wl_7 vdd gnd cell_6t
Xbit_r8_c248 bl_248 br_248 wl_8 vdd gnd cell_6t
Xbit_r9_c248 bl_248 br_248 wl_9 vdd gnd cell_6t
Xbit_r10_c248 bl_248 br_248 wl_10 vdd gnd cell_6t
Xbit_r11_c248 bl_248 br_248 wl_11 vdd gnd cell_6t
Xbit_r12_c248 bl_248 br_248 wl_12 vdd gnd cell_6t
Xbit_r13_c248 bl_248 br_248 wl_13 vdd gnd cell_6t
Xbit_r14_c248 bl_248 br_248 wl_14 vdd gnd cell_6t
Xbit_r15_c248 bl_248 br_248 wl_15 vdd gnd cell_6t
Xbit_r16_c248 bl_248 br_248 wl_16 vdd gnd cell_6t
Xbit_r17_c248 bl_248 br_248 wl_17 vdd gnd cell_6t
Xbit_r18_c248 bl_248 br_248 wl_18 vdd gnd cell_6t
Xbit_r19_c248 bl_248 br_248 wl_19 vdd gnd cell_6t
Xbit_r20_c248 bl_248 br_248 wl_20 vdd gnd cell_6t
Xbit_r21_c248 bl_248 br_248 wl_21 vdd gnd cell_6t
Xbit_r22_c248 bl_248 br_248 wl_22 vdd gnd cell_6t
Xbit_r23_c248 bl_248 br_248 wl_23 vdd gnd cell_6t
Xbit_r24_c248 bl_248 br_248 wl_24 vdd gnd cell_6t
Xbit_r25_c248 bl_248 br_248 wl_25 vdd gnd cell_6t
Xbit_r26_c248 bl_248 br_248 wl_26 vdd gnd cell_6t
Xbit_r27_c248 bl_248 br_248 wl_27 vdd gnd cell_6t
Xbit_r28_c248 bl_248 br_248 wl_28 vdd gnd cell_6t
Xbit_r29_c248 bl_248 br_248 wl_29 vdd gnd cell_6t
Xbit_r30_c248 bl_248 br_248 wl_30 vdd gnd cell_6t
Xbit_r31_c248 bl_248 br_248 wl_31 vdd gnd cell_6t
Xbit_r32_c248 bl_248 br_248 wl_32 vdd gnd cell_6t
Xbit_r33_c248 bl_248 br_248 wl_33 vdd gnd cell_6t
Xbit_r34_c248 bl_248 br_248 wl_34 vdd gnd cell_6t
Xbit_r35_c248 bl_248 br_248 wl_35 vdd gnd cell_6t
Xbit_r36_c248 bl_248 br_248 wl_36 vdd gnd cell_6t
Xbit_r37_c248 bl_248 br_248 wl_37 vdd gnd cell_6t
Xbit_r38_c248 bl_248 br_248 wl_38 vdd gnd cell_6t
Xbit_r39_c248 bl_248 br_248 wl_39 vdd gnd cell_6t
Xbit_r40_c248 bl_248 br_248 wl_40 vdd gnd cell_6t
Xbit_r41_c248 bl_248 br_248 wl_41 vdd gnd cell_6t
Xbit_r42_c248 bl_248 br_248 wl_42 vdd gnd cell_6t
Xbit_r43_c248 bl_248 br_248 wl_43 vdd gnd cell_6t
Xbit_r44_c248 bl_248 br_248 wl_44 vdd gnd cell_6t
Xbit_r45_c248 bl_248 br_248 wl_45 vdd gnd cell_6t
Xbit_r46_c248 bl_248 br_248 wl_46 vdd gnd cell_6t
Xbit_r47_c248 bl_248 br_248 wl_47 vdd gnd cell_6t
Xbit_r48_c248 bl_248 br_248 wl_48 vdd gnd cell_6t
Xbit_r49_c248 bl_248 br_248 wl_49 vdd gnd cell_6t
Xbit_r50_c248 bl_248 br_248 wl_50 vdd gnd cell_6t
Xbit_r51_c248 bl_248 br_248 wl_51 vdd gnd cell_6t
Xbit_r52_c248 bl_248 br_248 wl_52 vdd gnd cell_6t
Xbit_r53_c248 bl_248 br_248 wl_53 vdd gnd cell_6t
Xbit_r54_c248 bl_248 br_248 wl_54 vdd gnd cell_6t
Xbit_r55_c248 bl_248 br_248 wl_55 vdd gnd cell_6t
Xbit_r56_c248 bl_248 br_248 wl_56 vdd gnd cell_6t
Xbit_r57_c248 bl_248 br_248 wl_57 vdd gnd cell_6t
Xbit_r58_c248 bl_248 br_248 wl_58 vdd gnd cell_6t
Xbit_r59_c248 bl_248 br_248 wl_59 vdd gnd cell_6t
Xbit_r60_c248 bl_248 br_248 wl_60 vdd gnd cell_6t
Xbit_r61_c248 bl_248 br_248 wl_61 vdd gnd cell_6t
Xbit_r62_c248 bl_248 br_248 wl_62 vdd gnd cell_6t
Xbit_r63_c248 bl_248 br_248 wl_63 vdd gnd cell_6t
Xbit_r64_c248 bl_248 br_248 wl_64 vdd gnd cell_6t
Xbit_r65_c248 bl_248 br_248 wl_65 vdd gnd cell_6t
Xbit_r66_c248 bl_248 br_248 wl_66 vdd gnd cell_6t
Xbit_r67_c248 bl_248 br_248 wl_67 vdd gnd cell_6t
Xbit_r68_c248 bl_248 br_248 wl_68 vdd gnd cell_6t
Xbit_r69_c248 bl_248 br_248 wl_69 vdd gnd cell_6t
Xbit_r70_c248 bl_248 br_248 wl_70 vdd gnd cell_6t
Xbit_r71_c248 bl_248 br_248 wl_71 vdd gnd cell_6t
Xbit_r72_c248 bl_248 br_248 wl_72 vdd gnd cell_6t
Xbit_r73_c248 bl_248 br_248 wl_73 vdd gnd cell_6t
Xbit_r74_c248 bl_248 br_248 wl_74 vdd gnd cell_6t
Xbit_r75_c248 bl_248 br_248 wl_75 vdd gnd cell_6t
Xbit_r76_c248 bl_248 br_248 wl_76 vdd gnd cell_6t
Xbit_r77_c248 bl_248 br_248 wl_77 vdd gnd cell_6t
Xbit_r78_c248 bl_248 br_248 wl_78 vdd gnd cell_6t
Xbit_r79_c248 bl_248 br_248 wl_79 vdd gnd cell_6t
Xbit_r80_c248 bl_248 br_248 wl_80 vdd gnd cell_6t
Xbit_r81_c248 bl_248 br_248 wl_81 vdd gnd cell_6t
Xbit_r82_c248 bl_248 br_248 wl_82 vdd gnd cell_6t
Xbit_r83_c248 bl_248 br_248 wl_83 vdd gnd cell_6t
Xbit_r84_c248 bl_248 br_248 wl_84 vdd gnd cell_6t
Xbit_r85_c248 bl_248 br_248 wl_85 vdd gnd cell_6t
Xbit_r86_c248 bl_248 br_248 wl_86 vdd gnd cell_6t
Xbit_r87_c248 bl_248 br_248 wl_87 vdd gnd cell_6t
Xbit_r88_c248 bl_248 br_248 wl_88 vdd gnd cell_6t
Xbit_r89_c248 bl_248 br_248 wl_89 vdd gnd cell_6t
Xbit_r90_c248 bl_248 br_248 wl_90 vdd gnd cell_6t
Xbit_r91_c248 bl_248 br_248 wl_91 vdd gnd cell_6t
Xbit_r92_c248 bl_248 br_248 wl_92 vdd gnd cell_6t
Xbit_r93_c248 bl_248 br_248 wl_93 vdd gnd cell_6t
Xbit_r94_c248 bl_248 br_248 wl_94 vdd gnd cell_6t
Xbit_r95_c248 bl_248 br_248 wl_95 vdd gnd cell_6t
Xbit_r96_c248 bl_248 br_248 wl_96 vdd gnd cell_6t
Xbit_r97_c248 bl_248 br_248 wl_97 vdd gnd cell_6t
Xbit_r98_c248 bl_248 br_248 wl_98 vdd gnd cell_6t
Xbit_r99_c248 bl_248 br_248 wl_99 vdd gnd cell_6t
Xbit_r100_c248 bl_248 br_248 wl_100 vdd gnd cell_6t
Xbit_r101_c248 bl_248 br_248 wl_101 vdd gnd cell_6t
Xbit_r102_c248 bl_248 br_248 wl_102 vdd gnd cell_6t
Xbit_r103_c248 bl_248 br_248 wl_103 vdd gnd cell_6t
Xbit_r104_c248 bl_248 br_248 wl_104 vdd gnd cell_6t
Xbit_r105_c248 bl_248 br_248 wl_105 vdd gnd cell_6t
Xbit_r106_c248 bl_248 br_248 wl_106 vdd gnd cell_6t
Xbit_r107_c248 bl_248 br_248 wl_107 vdd gnd cell_6t
Xbit_r108_c248 bl_248 br_248 wl_108 vdd gnd cell_6t
Xbit_r109_c248 bl_248 br_248 wl_109 vdd gnd cell_6t
Xbit_r110_c248 bl_248 br_248 wl_110 vdd gnd cell_6t
Xbit_r111_c248 bl_248 br_248 wl_111 vdd gnd cell_6t
Xbit_r112_c248 bl_248 br_248 wl_112 vdd gnd cell_6t
Xbit_r113_c248 bl_248 br_248 wl_113 vdd gnd cell_6t
Xbit_r114_c248 bl_248 br_248 wl_114 vdd gnd cell_6t
Xbit_r115_c248 bl_248 br_248 wl_115 vdd gnd cell_6t
Xbit_r116_c248 bl_248 br_248 wl_116 vdd gnd cell_6t
Xbit_r117_c248 bl_248 br_248 wl_117 vdd gnd cell_6t
Xbit_r118_c248 bl_248 br_248 wl_118 vdd gnd cell_6t
Xbit_r119_c248 bl_248 br_248 wl_119 vdd gnd cell_6t
Xbit_r120_c248 bl_248 br_248 wl_120 vdd gnd cell_6t
Xbit_r121_c248 bl_248 br_248 wl_121 vdd gnd cell_6t
Xbit_r122_c248 bl_248 br_248 wl_122 vdd gnd cell_6t
Xbit_r123_c248 bl_248 br_248 wl_123 vdd gnd cell_6t
Xbit_r124_c248 bl_248 br_248 wl_124 vdd gnd cell_6t
Xbit_r125_c248 bl_248 br_248 wl_125 vdd gnd cell_6t
Xbit_r126_c248 bl_248 br_248 wl_126 vdd gnd cell_6t
Xbit_r127_c248 bl_248 br_248 wl_127 vdd gnd cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd cell_6t
Xbit_r1_c249 bl_249 br_249 wl_1 vdd gnd cell_6t
Xbit_r2_c249 bl_249 br_249 wl_2 vdd gnd cell_6t
Xbit_r3_c249 bl_249 br_249 wl_3 vdd gnd cell_6t
Xbit_r4_c249 bl_249 br_249 wl_4 vdd gnd cell_6t
Xbit_r5_c249 bl_249 br_249 wl_5 vdd gnd cell_6t
Xbit_r6_c249 bl_249 br_249 wl_6 vdd gnd cell_6t
Xbit_r7_c249 bl_249 br_249 wl_7 vdd gnd cell_6t
Xbit_r8_c249 bl_249 br_249 wl_8 vdd gnd cell_6t
Xbit_r9_c249 bl_249 br_249 wl_9 vdd gnd cell_6t
Xbit_r10_c249 bl_249 br_249 wl_10 vdd gnd cell_6t
Xbit_r11_c249 bl_249 br_249 wl_11 vdd gnd cell_6t
Xbit_r12_c249 bl_249 br_249 wl_12 vdd gnd cell_6t
Xbit_r13_c249 bl_249 br_249 wl_13 vdd gnd cell_6t
Xbit_r14_c249 bl_249 br_249 wl_14 vdd gnd cell_6t
Xbit_r15_c249 bl_249 br_249 wl_15 vdd gnd cell_6t
Xbit_r16_c249 bl_249 br_249 wl_16 vdd gnd cell_6t
Xbit_r17_c249 bl_249 br_249 wl_17 vdd gnd cell_6t
Xbit_r18_c249 bl_249 br_249 wl_18 vdd gnd cell_6t
Xbit_r19_c249 bl_249 br_249 wl_19 vdd gnd cell_6t
Xbit_r20_c249 bl_249 br_249 wl_20 vdd gnd cell_6t
Xbit_r21_c249 bl_249 br_249 wl_21 vdd gnd cell_6t
Xbit_r22_c249 bl_249 br_249 wl_22 vdd gnd cell_6t
Xbit_r23_c249 bl_249 br_249 wl_23 vdd gnd cell_6t
Xbit_r24_c249 bl_249 br_249 wl_24 vdd gnd cell_6t
Xbit_r25_c249 bl_249 br_249 wl_25 vdd gnd cell_6t
Xbit_r26_c249 bl_249 br_249 wl_26 vdd gnd cell_6t
Xbit_r27_c249 bl_249 br_249 wl_27 vdd gnd cell_6t
Xbit_r28_c249 bl_249 br_249 wl_28 vdd gnd cell_6t
Xbit_r29_c249 bl_249 br_249 wl_29 vdd gnd cell_6t
Xbit_r30_c249 bl_249 br_249 wl_30 vdd gnd cell_6t
Xbit_r31_c249 bl_249 br_249 wl_31 vdd gnd cell_6t
Xbit_r32_c249 bl_249 br_249 wl_32 vdd gnd cell_6t
Xbit_r33_c249 bl_249 br_249 wl_33 vdd gnd cell_6t
Xbit_r34_c249 bl_249 br_249 wl_34 vdd gnd cell_6t
Xbit_r35_c249 bl_249 br_249 wl_35 vdd gnd cell_6t
Xbit_r36_c249 bl_249 br_249 wl_36 vdd gnd cell_6t
Xbit_r37_c249 bl_249 br_249 wl_37 vdd gnd cell_6t
Xbit_r38_c249 bl_249 br_249 wl_38 vdd gnd cell_6t
Xbit_r39_c249 bl_249 br_249 wl_39 vdd gnd cell_6t
Xbit_r40_c249 bl_249 br_249 wl_40 vdd gnd cell_6t
Xbit_r41_c249 bl_249 br_249 wl_41 vdd gnd cell_6t
Xbit_r42_c249 bl_249 br_249 wl_42 vdd gnd cell_6t
Xbit_r43_c249 bl_249 br_249 wl_43 vdd gnd cell_6t
Xbit_r44_c249 bl_249 br_249 wl_44 vdd gnd cell_6t
Xbit_r45_c249 bl_249 br_249 wl_45 vdd gnd cell_6t
Xbit_r46_c249 bl_249 br_249 wl_46 vdd gnd cell_6t
Xbit_r47_c249 bl_249 br_249 wl_47 vdd gnd cell_6t
Xbit_r48_c249 bl_249 br_249 wl_48 vdd gnd cell_6t
Xbit_r49_c249 bl_249 br_249 wl_49 vdd gnd cell_6t
Xbit_r50_c249 bl_249 br_249 wl_50 vdd gnd cell_6t
Xbit_r51_c249 bl_249 br_249 wl_51 vdd gnd cell_6t
Xbit_r52_c249 bl_249 br_249 wl_52 vdd gnd cell_6t
Xbit_r53_c249 bl_249 br_249 wl_53 vdd gnd cell_6t
Xbit_r54_c249 bl_249 br_249 wl_54 vdd gnd cell_6t
Xbit_r55_c249 bl_249 br_249 wl_55 vdd gnd cell_6t
Xbit_r56_c249 bl_249 br_249 wl_56 vdd gnd cell_6t
Xbit_r57_c249 bl_249 br_249 wl_57 vdd gnd cell_6t
Xbit_r58_c249 bl_249 br_249 wl_58 vdd gnd cell_6t
Xbit_r59_c249 bl_249 br_249 wl_59 vdd gnd cell_6t
Xbit_r60_c249 bl_249 br_249 wl_60 vdd gnd cell_6t
Xbit_r61_c249 bl_249 br_249 wl_61 vdd gnd cell_6t
Xbit_r62_c249 bl_249 br_249 wl_62 vdd gnd cell_6t
Xbit_r63_c249 bl_249 br_249 wl_63 vdd gnd cell_6t
Xbit_r64_c249 bl_249 br_249 wl_64 vdd gnd cell_6t
Xbit_r65_c249 bl_249 br_249 wl_65 vdd gnd cell_6t
Xbit_r66_c249 bl_249 br_249 wl_66 vdd gnd cell_6t
Xbit_r67_c249 bl_249 br_249 wl_67 vdd gnd cell_6t
Xbit_r68_c249 bl_249 br_249 wl_68 vdd gnd cell_6t
Xbit_r69_c249 bl_249 br_249 wl_69 vdd gnd cell_6t
Xbit_r70_c249 bl_249 br_249 wl_70 vdd gnd cell_6t
Xbit_r71_c249 bl_249 br_249 wl_71 vdd gnd cell_6t
Xbit_r72_c249 bl_249 br_249 wl_72 vdd gnd cell_6t
Xbit_r73_c249 bl_249 br_249 wl_73 vdd gnd cell_6t
Xbit_r74_c249 bl_249 br_249 wl_74 vdd gnd cell_6t
Xbit_r75_c249 bl_249 br_249 wl_75 vdd gnd cell_6t
Xbit_r76_c249 bl_249 br_249 wl_76 vdd gnd cell_6t
Xbit_r77_c249 bl_249 br_249 wl_77 vdd gnd cell_6t
Xbit_r78_c249 bl_249 br_249 wl_78 vdd gnd cell_6t
Xbit_r79_c249 bl_249 br_249 wl_79 vdd gnd cell_6t
Xbit_r80_c249 bl_249 br_249 wl_80 vdd gnd cell_6t
Xbit_r81_c249 bl_249 br_249 wl_81 vdd gnd cell_6t
Xbit_r82_c249 bl_249 br_249 wl_82 vdd gnd cell_6t
Xbit_r83_c249 bl_249 br_249 wl_83 vdd gnd cell_6t
Xbit_r84_c249 bl_249 br_249 wl_84 vdd gnd cell_6t
Xbit_r85_c249 bl_249 br_249 wl_85 vdd gnd cell_6t
Xbit_r86_c249 bl_249 br_249 wl_86 vdd gnd cell_6t
Xbit_r87_c249 bl_249 br_249 wl_87 vdd gnd cell_6t
Xbit_r88_c249 bl_249 br_249 wl_88 vdd gnd cell_6t
Xbit_r89_c249 bl_249 br_249 wl_89 vdd gnd cell_6t
Xbit_r90_c249 bl_249 br_249 wl_90 vdd gnd cell_6t
Xbit_r91_c249 bl_249 br_249 wl_91 vdd gnd cell_6t
Xbit_r92_c249 bl_249 br_249 wl_92 vdd gnd cell_6t
Xbit_r93_c249 bl_249 br_249 wl_93 vdd gnd cell_6t
Xbit_r94_c249 bl_249 br_249 wl_94 vdd gnd cell_6t
Xbit_r95_c249 bl_249 br_249 wl_95 vdd gnd cell_6t
Xbit_r96_c249 bl_249 br_249 wl_96 vdd gnd cell_6t
Xbit_r97_c249 bl_249 br_249 wl_97 vdd gnd cell_6t
Xbit_r98_c249 bl_249 br_249 wl_98 vdd gnd cell_6t
Xbit_r99_c249 bl_249 br_249 wl_99 vdd gnd cell_6t
Xbit_r100_c249 bl_249 br_249 wl_100 vdd gnd cell_6t
Xbit_r101_c249 bl_249 br_249 wl_101 vdd gnd cell_6t
Xbit_r102_c249 bl_249 br_249 wl_102 vdd gnd cell_6t
Xbit_r103_c249 bl_249 br_249 wl_103 vdd gnd cell_6t
Xbit_r104_c249 bl_249 br_249 wl_104 vdd gnd cell_6t
Xbit_r105_c249 bl_249 br_249 wl_105 vdd gnd cell_6t
Xbit_r106_c249 bl_249 br_249 wl_106 vdd gnd cell_6t
Xbit_r107_c249 bl_249 br_249 wl_107 vdd gnd cell_6t
Xbit_r108_c249 bl_249 br_249 wl_108 vdd gnd cell_6t
Xbit_r109_c249 bl_249 br_249 wl_109 vdd gnd cell_6t
Xbit_r110_c249 bl_249 br_249 wl_110 vdd gnd cell_6t
Xbit_r111_c249 bl_249 br_249 wl_111 vdd gnd cell_6t
Xbit_r112_c249 bl_249 br_249 wl_112 vdd gnd cell_6t
Xbit_r113_c249 bl_249 br_249 wl_113 vdd gnd cell_6t
Xbit_r114_c249 bl_249 br_249 wl_114 vdd gnd cell_6t
Xbit_r115_c249 bl_249 br_249 wl_115 vdd gnd cell_6t
Xbit_r116_c249 bl_249 br_249 wl_116 vdd gnd cell_6t
Xbit_r117_c249 bl_249 br_249 wl_117 vdd gnd cell_6t
Xbit_r118_c249 bl_249 br_249 wl_118 vdd gnd cell_6t
Xbit_r119_c249 bl_249 br_249 wl_119 vdd gnd cell_6t
Xbit_r120_c249 bl_249 br_249 wl_120 vdd gnd cell_6t
Xbit_r121_c249 bl_249 br_249 wl_121 vdd gnd cell_6t
Xbit_r122_c249 bl_249 br_249 wl_122 vdd gnd cell_6t
Xbit_r123_c249 bl_249 br_249 wl_123 vdd gnd cell_6t
Xbit_r124_c249 bl_249 br_249 wl_124 vdd gnd cell_6t
Xbit_r125_c249 bl_249 br_249 wl_125 vdd gnd cell_6t
Xbit_r126_c249 bl_249 br_249 wl_126 vdd gnd cell_6t
Xbit_r127_c249 bl_249 br_249 wl_127 vdd gnd cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd cell_6t
Xbit_r1_c250 bl_250 br_250 wl_1 vdd gnd cell_6t
Xbit_r2_c250 bl_250 br_250 wl_2 vdd gnd cell_6t
Xbit_r3_c250 bl_250 br_250 wl_3 vdd gnd cell_6t
Xbit_r4_c250 bl_250 br_250 wl_4 vdd gnd cell_6t
Xbit_r5_c250 bl_250 br_250 wl_5 vdd gnd cell_6t
Xbit_r6_c250 bl_250 br_250 wl_6 vdd gnd cell_6t
Xbit_r7_c250 bl_250 br_250 wl_7 vdd gnd cell_6t
Xbit_r8_c250 bl_250 br_250 wl_8 vdd gnd cell_6t
Xbit_r9_c250 bl_250 br_250 wl_9 vdd gnd cell_6t
Xbit_r10_c250 bl_250 br_250 wl_10 vdd gnd cell_6t
Xbit_r11_c250 bl_250 br_250 wl_11 vdd gnd cell_6t
Xbit_r12_c250 bl_250 br_250 wl_12 vdd gnd cell_6t
Xbit_r13_c250 bl_250 br_250 wl_13 vdd gnd cell_6t
Xbit_r14_c250 bl_250 br_250 wl_14 vdd gnd cell_6t
Xbit_r15_c250 bl_250 br_250 wl_15 vdd gnd cell_6t
Xbit_r16_c250 bl_250 br_250 wl_16 vdd gnd cell_6t
Xbit_r17_c250 bl_250 br_250 wl_17 vdd gnd cell_6t
Xbit_r18_c250 bl_250 br_250 wl_18 vdd gnd cell_6t
Xbit_r19_c250 bl_250 br_250 wl_19 vdd gnd cell_6t
Xbit_r20_c250 bl_250 br_250 wl_20 vdd gnd cell_6t
Xbit_r21_c250 bl_250 br_250 wl_21 vdd gnd cell_6t
Xbit_r22_c250 bl_250 br_250 wl_22 vdd gnd cell_6t
Xbit_r23_c250 bl_250 br_250 wl_23 vdd gnd cell_6t
Xbit_r24_c250 bl_250 br_250 wl_24 vdd gnd cell_6t
Xbit_r25_c250 bl_250 br_250 wl_25 vdd gnd cell_6t
Xbit_r26_c250 bl_250 br_250 wl_26 vdd gnd cell_6t
Xbit_r27_c250 bl_250 br_250 wl_27 vdd gnd cell_6t
Xbit_r28_c250 bl_250 br_250 wl_28 vdd gnd cell_6t
Xbit_r29_c250 bl_250 br_250 wl_29 vdd gnd cell_6t
Xbit_r30_c250 bl_250 br_250 wl_30 vdd gnd cell_6t
Xbit_r31_c250 bl_250 br_250 wl_31 vdd gnd cell_6t
Xbit_r32_c250 bl_250 br_250 wl_32 vdd gnd cell_6t
Xbit_r33_c250 bl_250 br_250 wl_33 vdd gnd cell_6t
Xbit_r34_c250 bl_250 br_250 wl_34 vdd gnd cell_6t
Xbit_r35_c250 bl_250 br_250 wl_35 vdd gnd cell_6t
Xbit_r36_c250 bl_250 br_250 wl_36 vdd gnd cell_6t
Xbit_r37_c250 bl_250 br_250 wl_37 vdd gnd cell_6t
Xbit_r38_c250 bl_250 br_250 wl_38 vdd gnd cell_6t
Xbit_r39_c250 bl_250 br_250 wl_39 vdd gnd cell_6t
Xbit_r40_c250 bl_250 br_250 wl_40 vdd gnd cell_6t
Xbit_r41_c250 bl_250 br_250 wl_41 vdd gnd cell_6t
Xbit_r42_c250 bl_250 br_250 wl_42 vdd gnd cell_6t
Xbit_r43_c250 bl_250 br_250 wl_43 vdd gnd cell_6t
Xbit_r44_c250 bl_250 br_250 wl_44 vdd gnd cell_6t
Xbit_r45_c250 bl_250 br_250 wl_45 vdd gnd cell_6t
Xbit_r46_c250 bl_250 br_250 wl_46 vdd gnd cell_6t
Xbit_r47_c250 bl_250 br_250 wl_47 vdd gnd cell_6t
Xbit_r48_c250 bl_250 br_250 wl_48 vdd gnd cell_6t
Xbit_r49_c250 bl_250 br_250 wl_49 vdd gnd cell_6t
Xbit_r50_c250 bl_250 br_250 wl_50 vdd gnd cell_6t
Xbit_r51_c250 bl_250 br_250 wl_51 vdd gnd cell_6t
Xbit_r52_c250 bl_250 br_250 wl_52 vdd gnd cell_6t
Xbit_r53_c250 bl_250 br_250 wl_53 vdd gnd cell_6t
Xbit_r54_c250 bl_250 br_250 wl_54 vdd gnd cell_6t
Xbit_r55_c250 bl_250 br_250 wl_55 vdd gnd cell_6t
Xbit_r56_c250 bl_250 br_250 wl_56 vdd gnd cell_6t
Xbit_r57_c250 bl_250 br_250 wl_57 vdd gnd cell_6t
Xbit_r58_c250 bl_250 br_250 wl_58 vdd gnd cell_6t
Xbit_r59_c250 bl_250 br_250 wl_59 vdd gnd cell_6t
Xbit_r60_c250 bl_250 br_250 wl_60 vdd gnd cell_6t
Xbit_r61_c250 bl_250 br_250 wl_61 vdd gnd cell_6t
Xbit_r62_c250 bl_250 br_250 wl_62 vdd gnd cell_6t
Xbit_r63_c250 bl_250 br_250 wl_63 vdd gnd cell_6t
Xbit_r64_c250 bl_250 br_250 wl_64 vdd gnd cell_6t
Xbit_r65_c250 bl_250 br_250 wl_65 vdd gnd cell_6t
Xbit_r66_c250 bl_250 br_250 wl_66 vdd gnd cell_6t
Xbit_r67_c250 bl_250 br_250 wl_67 vdd gnd cell_6t
Xbit_r68_c250 bl_250 br_250 wl_68 vdd gnd cell_6t
Xbit_r69_c250 bl_250 br_250 wl_69 vdd gnd cell_6t
Xbit_r70_c250 bl_250 br_250 wl_70 vdd gnd cell_6t
Xbit_r71_c250 bl_250 br_250 wl_71 vdd gnd cell_6t
Xbit_r72_c250 bl_250 br_250 wl_72 vdd gnd cell_6t
Xbit_r73_c250 bl_250 br_250 wl_73 vdd gnd cell_6t
Xbit_r74_c250 bl_250 br_250 wl_74 vdd gnd cell_6t
Xbit_r75_c250 bl_250 br_250 wl_75 vdd gnd cell_6t
Xbit_r76_c250 bl_250 br_250 wl_76 vdd gnd cell_6t
Xbit_r77_c250 bl_250 br_250 wl_77 vdd gnd cell_6t
Xbit_r78_c250 bl_250 br_250 wl_78 vdd gnd cell_6t
Xbit_r79_c250 bl_250 br_250 wl_79 vdd gnd cell_6t
Xbit_r80_c250 bl_250 br_250 wl_80 vdd gnd cell_6t
Xbit_r81_c250 bl_250 br_250 wl_81 vdd gnd cell_6t
Xbit_r82_c250 bl_250 br_250 wl_82 vdd gnd cell_6t
Xbit_r83_c250 bl_250 br_250 wl_83 vdd gnd cell_6t
Xbit_r84_c250 bl_250 br_250 wl_84 vdd gnd cell_6t
Xbit_r85_c250 bl_250 br_250 wl_85 vdd gnd cell_6t
Xbit_r86_c250 bl_250 br_250 wl_86 vdd gnd cell_6t
Xbit_r87_c250 bl_250 br_250 wl_87 vdd gnd cell_6t
Xbit_r88_c250 bl_250 br_250 wl_88 vdd gnd cell_6t
Xbit_r89_c250 bl_250 br_250 wl_89 vdd gnd cell_6t
Xbit_r90_c250 bl_250 br_250 wl_90 vdd gnd cell_6t
Xbit_r91_c250 bl_250 br_250 wl_91 vdd gnd cell_6t
Xbit_r92_c250 bl_250 br_250 wl_92 vdd gnd cell_6t
Xbit_r93_c250 bl_250 br_250 wl_93 vdd gnd cell_6t
Xbit_r94_c250 bl_250 br_250 wl_94 vdd gnd cell_6t
Xbit_r95_c250 bl_250 br_250 wl_95 vdd gnd cell_6t
Xbit_r96_c250 bl_250 br_250 wl_96 vdd gnd cell_6t
Xbit_r97_c250 bl_250 br_250 wl_97 vdd gnd cell_6t
Xbit_r98_c250 bl_250 br_250 wl_98 vdd gnd cell_6t
Xbit_r99_c250 bl_250 br_250 wl_99 vdd gnd cell_6t
Xbit_r100_c250 bl_250 br_250 wl_100 vdd gnd cell_6t
Xbit_r101_c250 bl_250 br_250 wl_101 vdd gnd cell_6t
Xbit_r102_c250 bl_250 br_250 wl_102 vdd gnd cell_6t
Xbit_r103_c250 bl_250 br_250 wl_103 vdd gnd cell_6t
Xbit_r104_c250 bl_250 br_250 wl_104 vdd gnd cell_6t
Xbit_r105_c250 bl_250 br_250 wl_105 vdd gnd cell_6t
Xbit_r106_c250 bl_250 br_250 wl_106 vdd gnd cell_6t
Xbit_r107_c250 bl_250 br_250 wl_107 vdd gnd cell_6t
Xbit_r108_c250 bl_250 br_250 wl_108 vdd gnd cell_6t
Xbit_r109_c250 bl_250 br_250 wl_109 vdd gnd cell_6t
Xbit_r110_c250 bl_250 br_250 wl_110 vdd gnd cell_6t
Xbit_r111_c250 bl_250 br_250 wl_111 vdd gnd cell_6t
Xbit_r112_c250 bl_250 br_250 wl_112 vdd gnd cell_6t
Xbit_r113_c250 bl_250 br_250 wl_113 vdd gnd cell_6t
Xbit_r114_c250 bl_250 br_250 wl_114 vdd gnd cell_6t
Xbit_r115_c250 bl_250 br_250 wl_115 vdd gnd cell_6t
Xbit_r116_c250 bl_250 br_250 wl_116 vdd gnd cell_6t
Xbit_r117_c250 bl_250 br_250 wl_117 vdd gnd cell_6t
Xbit_r118_c250 bl_250 br_250 wl_118 vdd gnd cell_6t
Xbit_r119_c250 bl_250 br_250 wl_119 vdd gnd cell_6t
Xbit_r120_c250 bl_250 br_250 wl_120 vdd gnd cell_6t
Xbit_r121_c250 bl_250 br_250 wl_121 vdd gnd cell_6t
Xbit_r122_c250 bl_250 br_250 wl_122 vdd gnd cell_6t
Xbit_r123_c250 bl_250 br_250 wl_123 vdd gnd cell_6t
Xbit_r124_c250 bl_250 br_250 wl_124 vdd gnd cell_6t
Xbit_r125_c250 bl_250 br_250 wl_125 vdd gnd cell_6t
Xbit_r126_c250 bl_250 br_250 wl_126 vdd gnd cell_6t
Xbit_r127_c250 bl_250 br_250 wl_127 vdd gnd cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd cell_6t
Xbit_r1_c251 bl_251 br_251 wl_1 vdd gnd cell_6t
Xbit_r2_c251 bl_251 br_251 wl_2 vdd gnd cell_6t
Xbit_r3_c251 bl_251 br_251 wl_3 vdd gnd cell_6t
Xbit_r4_c251 bl_251 br_251 wl_4 vdd gnd cell_6t
Xbit_r5_c251 bl_251 br_251 wl_5 vdd gnd cell_6t
Xbit_r6_c251 bl_251 br_251 wl_6 vdd gnd cell_6t
Xbit_r7_c251 bl_251 br_251 wl_7 vdd gnd cell_6t
Xbit_r8_c251 bl_251 br_251 wl_8 vdd gnd cell_6t
Xbit_r9_c251 bl_251 br_251 wl_9 vdd gnd cell_6t
Xbit_r10_c251 bl_251 br_251 wl_10 vdd gnd cell_6t
Xbit_r11_c251 bl_251 br_251 wl_11 vdd gnd cell_6t
Xbit_r12_c251 bl_251 br_251 wl_12 vdd gnd cell_6t
Xbit_r13_c251 bl_251 br_251 wl_13 vdd gnd cell_6t
Xbit_r14_c251 bl_251 br_251 wl_14 vdd gnd cell_6t
Xbit_r15_c251 bl_251 br_251 wl_15 vdd gnd cell_6t
Xbit_r16_c251 bl_251 br_251 wl_16 vdd gnd cell_6t
Xbit_r17_c251 bl_251 br_251 wl_17 vdd gnd cell_6t
Xbit_r18_c251 bl_251 br_251 wl_18 vdd gnd cell_6t
Xbit_r19_c251 bl_251 br_251 wl_19 vdd gnd cell_6t
Xbit_r20_c251 bl_251 br_251 wl_20 vdd gnd cell_6t
Xbit_r21_c251 bl_251 br_251 wl_21 vdd gnd cell_6t
Xbit_r22_c251 bl_251 br_251 wl_22 vdd gnd cell_6t
Xbit_r23_c251 bl_251 br_251 wl_23 vdd gnd cell_6t
Xbit_r24_c251 bl_251 br_251 wl_24 vdd gnd cell_6t
Xbit_r25_c251 bl_251 br_251 wl_25 vdd gnd cell_6t
Xbit_r26_c251 bl_251 br_251 wl_26 vdd gnd cell_6t
Xbit_r27_c251 bl_251 br_251 wl_27 vdd gnd cell_6t
Xbit_r28_c251 bl_251 br_251 wl_28 vdd gnd cell_6t
Xbit_r29_c251 bl_251 br_251 wl_29 vdd gnd cell_6t
Xbit_r30_c251 bl_251 br_251 wl_30 vdd gnd cell_6t
Xbit_r31_c251 bl_251 br_251 wl_31 vdd gnd cell_6t
Xbit_r32_c251 bl_251 br_251 wl_32 vdd gnd cell_6t
Xbit_r33_c251 bl_251 br_251 wl_33 vdd gnd cell_6t
Xbit_r34_c251 bl_251 br_251 wl_34 vdd gnd cell_6t
Xbit_r35_c251 bl_251 br_251 wl_35 vdd gnd cell_6t
Xbit_r36_c251 bl_251 br_251 wl_36 vdd gnd cell_6t
Xbit_r37_c251 bl_251 br_251 wl_37 vdd gnd cell_6t
Xbit_r38_c251 bl_251 br_251 wl_38 vdd gnd cell_6t
Xbit_r39_c251 bl_251 br_251 wl_39 vdd gnd cell_6t
Xbit_r40_c251 bl_251 br_251 wl_40 vdd gnd cell_6t
Xbit_r41_c251 bl_251 br_251 wl_41 vdd gnd cell_6t
Xbit_r42_c251 bl_251 br_251 wl_42 vdd gnd cell_6t
Xbit_r43_c251 bl_251 br_251 wl_43 vdd gnd cell_6t
Xbit_r44_c251 bl_251 br_251 wl_44 vdd gnd cell_6t
Xbit_r45_c251 bl_251 br_251 wl_45 vdd gnd cell_6t
Xbit_r46_c251 bl_251 br_251 wl_46 vdd gnd cell_6t
Xbit_r47_c251 bl_251 br_251 wl_47 vdd gnd cell_6t
Xbit_r48_c251 bl_251 br_251 wl_48 vdd gnd cell_6t
Xbit_r49_c251 bl_251 br_251 wl_49 vdd gnd cell_6t
Xbit_r50_c251 bl_251 br_251 wl_50 vdd gnd cell_6t
Xbit_r51_c251 bl_251 br_251 wl_51 vdd gnd cell_6t
Xbit_r52_c251 bl_251 br_251 wl_52 vdd gnd cell_6t
Xbit_r53_c251 bl_251 br_251 wl_53 vdd gnd cell_6t
Xbit_r54_c251 bl_251 br_251 wl_54 vdd gnd cell_6t
Xbit_r55_c251 bl_251 br_251 wl_55 vdd gnd cell_6t
Xbit_r56_c251 bl_251 br_251 wl_56 vdd gnd cell_6t
Xbit_r57_c251 bl_251 br_251 wl_57 vdd gnd cell_6t
Xbit_r58_c251 bl_251 br_251 wl_58 vdd gnd cell_6t
Xbit_r59_c251 bl_251 br_251 wl_59 vdd gnd cell_6t
Xbit_r60_c251 bl_251 br_251 wl_60 vdd gnd cell_6t
Xbit_r61_c251 bl_251 br_251 wl_61 vdd gnd cell_6t
Xbit_r62_c251 bl_251 br_251 wl_62 vdd gnd cell_6t
Xbit_r63_c251 bl_251 br_251 wl_63 vdd gnd cell_6t
Xbit_r64_c251 bl_251 br_251 wl_64 vdd gnd cell_6t
Xbit_r65_c251 bl_251 br_251 wl_65 vdd gnd cell_6t
Xbit_r66_c251 bl_251 br_251 wl_66 vdd gnd cell_6t
Xbit_r67_c251 bl_251 br_251 wl_67 vdd gnd cell_6t
Xbit_r68_c251 bl_251 br_251 wl_68 vdd gnd cell_6t
Xbit_r69_c251 bl_251 br_251 wl_69 vdd gnd cell_6t
Xbit_r70_c251 bl_251 br_251 wl_70 vdd gnd cell_6t
Xbit_r71_c251 bl_251 br_251 wl_71 vdd gnd cell_6t
Xbit_r72_c251 bl_251 br_251 wl_72 vdd gnd cell_6t
Xbit_r73_c251 bl_251 br_251 wl_73 vdd gnd cell_6t
Xbit_r74_c251 bl_251 br_251 wl_74 vdd gnd cell_6t
Xbit_r75_c251 bl_251 br_251 wl_75 vdd gnd cell_6t
Xbit_r76_c251 bl_251 br_251 wl_76 vdd gnd cell_6t
Xbit_r77_c251 bl_251 br_251 wl_77 vdd gnd cell_6t
Xbit_r78_c251 bl_251 br_251 wl_78 vdd gnd cell_6t
Xbit_r79_c251 bl_251 br_251 wl_79 vdd gnd cell_6t
Xbit_r80_c251 bl_251 br_251 wl_80 vdd gnd cell_6t
Xbit_r81_c251 bl_251 br_251 wl_81 vdd gnd cell_6t
Xbit_r82_c251 bl_251 br_251 wl_82 vdd gnd cell_6t
Xbit_r83_c251 bl_251 br_251 wl_83 vdd gnd cell_6t
Xbit_r84_c251 bl_251 br_251 wl_84 vdd gnd cell_6t
Xbit_r85_c251 bl_251 br_251 wl_85 vdd gnd cell_6t
Xbit_r86_c251 bl_251 br_251 wl_86 vdd gnd cell_6t
Xbit_r87_c251 bl_251 br_251 wl_87 vdd gnd cell_6t
Xbit_r88_c251 bl_251 br_251 wl_88 vdd gnd cell_6t
Xbit_r89_c251 bl_251 br_251 wl_89 vdd gnd cell_6t
Xbit_r90_c251 bl_251 br_251 wl_90 vdd gnd cell_6t
Xbit_r91_c251 bl_251 br_251 wl_91 vdd gnd cell_6t
Xbit_r92_c251 bl_251 br_251 wl_92 vdd gnd cell_6t
Xbit_r93_c251 bl_251 br_251 wl_93 vdd gnd cell_6t
Xbit_r94_c251 bl_251 br_251 wl_94 vdd gnd cell_6t
Xbit_r95_c251 bl_251 br_251 wl_95 vdd gnd cell_6t
Xbit_r96_c251 bl_251 br_251 wl_96 vdd gnd cell_6t
Xbit_r97_c251 bl_251 br_251 wl_97 vdd gnd cell_6t
Xbit_r98_c251 bl_251 br_251 wl_98 vdd gnd cell_6t
Xbit_r99_c251 bl_251 br_251 wl_99 vdd gnd cell_6t
Xbit_r100_c251 bl_251 br_251 wl_100 vdd gnd cell_6t
Xbit_r101_c251 bl_251 br_251 wl_101 vdd gnd cell_6t
Xbit_r102_c251 bl_251 br_251 wl_102 vdd gnd cell_6t
Xbit_r103_c251 bl_251 br_251 wl_103 vdd gnd cell_6t
Xbit_r104_c251 bl_251 br_251 wl_104 vdd gnd cell_6t
Xbit_r105_c251 bl_251 br_251 wl_105 vdd gnd cell_6t
Xbit_r106_c251 bl_251 br_251 wl_106 vdd gnd cell_6t
Xbit_r107_c251 bl_251 br_251 wl_107 vdd gnd cell_6t
Xbit_r108_c251 bl_251 br_251 wl_108 vdd gnd cell_6t
Xbit_r109_c251 bl_251 br_251 wl_109 vdd gnd cell_6t
Xbit_r110_c251 bl_251 br_251 wl_110 vdd gnd cell_6t
Xbit_r111_c251 bl_251 br_251 wl_111 vdd gnd cell_6t
Xbit_r112_c251 bl_251 br_251 wl_112 vdd gnd cell_6t
Xbit_r113_c251 bl_251 br_251 wl_113 vdd gnd cell_6t
Xbit_r114_c251 bl_251 br_251 wl_114 vdd gnd cell_6t
Xbit_r115_c251 bl_251 br_251 wl_115 vdd gnd cell_6t
Xbit_r116_c251 bl_251 br_251 wl_116 vdd gnd cell_6t
Xbit_r117_c251 bl_251 br_251 wl_117 vdd gnd cell_6t
Xbit_r118_c251 bl_251 br_251 wl_118 vdd gnd cell_6t
Xbit_r119_c251 bl_251 br_251 wl_119 vdd gnd cell_6t
Xbit_r120_c251 bl_251 br_251 wl_120 vdd gnd cell_6t
Xbit_r121_c251 bl_251 br_251 wl_121 vdd gnd cell_6t
Xbit_r122_c251 bl_251 br_251 wl_122 vdd gnd cell_6t
Xbit_r123_c251 bl_251 br_251 wl_123 vdd gnd cell_6t
Xbit_r124_c251 bl_251 br_251 wl_124 vdd gnd cell_6t
Xbit_r125_c251 bl_251 br_251 wl_125 vdd gnd cell_6t
Xbit_r126_c251 bl_251 br_251 wl_126 vdd gnd cell_6t
Xbit_r127_c251 bl_251 br_251 wl_127 vdd gnd cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd cell_6t
Xbit_r1_c252 bl_252 br_252 wl_1 vdd gnd cell_6t
Xbit_r2_c252 bl_252 br_252 wl_2 vdd gnd cell_6t
Xbit_r3_c252 bl_252 br_252 wl_3 vdd gnd cell_6t
Xbit_r4_c252 bl_252 br_252 wl_4 vdd gnd cell_6t
Xbit_r5_c252 bl_252 br_252 wl_5 vdd gnd cell_6t
Xbit_r6_c252 bl_252 br_252 wl_6 vdd gnd cell_6t
Xbit_r7_c252 bl_252 br_252 wl_7 vdd gnd cell_6t
Xbit_r8_c252 bl_252 br_252 wl_8 vdd gnd cell_6t
Xbit_r9_c252 bl_252 br_252 wl_9 vdd gnd cell_6t
Xbit_r10_c252 bl_252 br_252 wl_10 vdd gnd cell_6t
Xbit_r11_c252 bl_252 br_252 wl_11 vdd gnd cell_6t
Xbit_r12_c252 bl_252 br_252 wl_12 vdd gnd cell_6t
Xbit_r13_c252 bl_252 br_252 wl_13 vdd gnd cell_6t
Xbit_r14_c252 bl_252 br_252 wl_14 vdd gnd cell_6t
Xbit_r15_c252 bl_252 br_252 wl_15 vdd gnd cell_6t
Xbit_r16_c252 bl_252 br_252 wl_16 vdd gnd cell_6t
Xbit_r17_c252 bl_252 br_252 wl_17 vdd gnd cell_6t
Xbit_r18_c252 bl_252 br_252 wl_18 vdd gnd cell_6t
Xbit_r19_c252 bl_252 br_252 wl_19 vdd gnd cell_6t
Xbit_r20_c252 bl_252 br_252 wl_20 vdd gnd cell_6t
Xbit_r21_c252 bl_252 br_252 wl_21 vdd gnd cell_6t
Xbit_r22_c252 bl_252 br_252 wl_22 vdd gnd cell_6t
Xbit_r23_c252 bl_252 br_252 wl_23 vdd gnd cell_6t
Xbit_r24_c252 bl_252 br_252 wl_24 vdd gnd cell_6t
Xbit_r25_c252 bl_252 br_252 wl_25 vdd gnd cell_6t
Xbit_r26_c252 bl_252 br_252 wl_26 vdd gnd cell_6t
Xbit_r27_c252 bl_252 br_252 wl_27 vdd gnd cell_6t
Xbit_r28_c252 bl_252 br_252 wl_28 vdd gnd cell_6t
Xbit_r29_c252 bl_252 br_252 wl_29 vdd gnd cell_6t
Xbit_r30_c252 bl_252 br_252 wl_30 vdd gnd cell_6t
Xbit_r31_c252 bl_252 br_252 wl_31 vdd gnd cell_6t
Xbit_r32_c252 bl_252 br_252 wl_32 vdd gnd cell_6t
Xbit_r33_c252 bl_252 br_252 wl_33 vdd gnd cell_6t
Xbit_r34_c252 bl_252 br_252 wl_34 vdd gnd cell_6t
Xbit_r35_c252 bl_252 br_252 wl_35 vdd gnd cell_6t
Xbit_r36_c252 bl_252 br_252 wl_36 vdd gnd cell_6t
Xbit_r37_c252 bl_252 br_252 wl_37 vdd gnd cell_6t
Xbit_r38_c252 bl_252 br_252 wl_38 vdd gnd cell_6t
Xbit_r39_c252 bl_252 br_252 wl_39 vdd gnd cell_6t
Xbit_r40_c252 bl_252 br_252 wl_40 vdd gnd cell_6t
Xbit_r41_c252 bl_252 br_252 wl_41 vdd gnd cell_6t
Xbit_r42_c252 bl_252 br_252 wl_42 vdd gnd cell_6t
Xbit_r43_c252 bl_252 br_252 wl_43 vdd gnd cell_6t
Xbit_r44_c252 bl_252 br_252 wl_44 vdd gnd cell_6t
Xbit_r45_c252 bl_252 br_252 wl_45 vdd gnd cell_6t
Xbit_r46_c252 bl_252 br_252 wl_46 vdd gnd cell_6t
Xbit_r47_c252 bl_252 br_252 wl_47 vdd gnd cell_6t
Xbit_r48_c252 bl_252 br_252 wl_48 vdd gnd cell_6t
Xbit_r49_c252 bl_252 br_252 wl_49 vdd gnd cell_6t
Xbit_r50_c252 bl_252 br_252 wl_50 vdd gnd cell_6t
Xbit_r51_c252 bl_252 br_252 wl_51 vdd gnd cell_6t
Xbit_r52_c252 bl_252 br_252 wl_52 vdd gnd cell_6t
Xbit_r53_c252 bl_252 br_252 wl_53 vdd gnd cell_6t
Xbit_r54_c252 bl_252 br_252 wl_54 vdd gnd cell_6t
Xbit_r55_c252 bl_252 br_252 wl_55 vdd gnd cell_6t
Xbit_r56_c252 bl_252 br_252 wl_56 vdd gnd cell_6t
Xbit_r57_c252 bl_252 br_252 wl_57 vdd gnd cell_6t
Xbit_r58_c252 bl_252 br_252 wl_58 vdd gnd cell_6t
Xbit_r59_c252 bl_252 br_252 wl_59 vdd gnd cell_6t
Xbit_r60_c252 bl_252 br_252 wl_60 vdd gnd cell_6t
Xbit_r61_c252 bl_252 br_252 wl_61 vdd gnd cell_6t
Xbit_r62_c252 bl_252 br_252 wl_62 vdd gnd cell_6t
Xbit_r63_c252 bl_252 br_252 wl_63 vdd gnd cell_6t
Xbit_r64_c252 bl_252 br_252 wl_64 vdd gnd cell_6t
Xbit_r65_c252 bl_252 br_252 wl_65 vdd gnd cell_6t
Xbit_r66_c252 bl_252 br_252 wl_66 vdd gnd cell_6t
Xbit_r67_c252 bl_252 br_252 wl_67 vdd gnd cell_6t
Xbit_r68_c252 bl_252 br_252 wl_68 vdd gnd cell_6t
Xbit_r69_c252 bl_252 br_252 wl_69 vdd gnd cell_6t
Xbit_r70_c252 bl_252 br_252 wl_70 vdd gnd cell_6t
Xbit_r71_c252 bl_252 br_252 wl_71 vdd gnd cell_6t
Xbit_r72_c252 bl_252 br_252 wl_72 vdd gnd cell_6t
Xbit_r73_c252 bl_252 br_252 wl_73 vdd gnd cell_6t
Xbit_r74_c252 bl_252 br_252 wl_74 vdd gnd cell_6t
Xbit_r75_c252 bl_252 br_252 wl_75 vdd gnd cell_6t
Xbit_r76_c252 bl_252 br_252 wl_76 vdd gnd cell_6t
Xbit_r77_c252 bl_252 br_252 wl_77 vdd gnd cell_6t
Xbit_r78_c252 bl_252 br_252 wl_78 vdd gnd cell_6t
Xbit_r79_c252 bl_252 br_252 wl_79 vdd gnd cell_6t
Xbit_r80_c252 bl_252 br_252 wl_80 vdd gnd cell_6t
Xbit_r81_c252 bl_252 br_252 wl_81 vdd gnd cell_6t
Xbit_r82_c252 bl_252 br_252 wl_82 vdd gnd cell_6t
Xbit_r83_c252 bl_252 br_252 wl_83 vdd gnd cell_6t
Xbit_r84_c252 bl_252 br_252 wl_84 vdd gnd cell_6t
Xbit_r85_c252 bl_252 br_252 wl_85 vdd gnd cell_6t
Xbit_r86_c252 bl_252 br_252 wl_86 vdd gnd cell_6t
Xbit_r87_c252 bl_252 br_252 wl_87 vdd gnd cell_6t
Xbit_r88_c252 bl_252 br_252 wl_88 vdd gnd cell_6t
Xbit_r89_c252 bl_252 br_252 wl_89 vdd gnd cell_6t
Xbit_r90_c252 bl_252 br_252 wl_90 vdd gnd cell_6t
Xbit_r91_c252 bl_252 br_252 wl_91 vdd gnd cell_6t
Xbit_r92_c252 bl_252 br_252 wl_92 vdd gnd cell_6t
Xbit_r93_c252 bl_252 br_252 wl_93 vdd gnd cell_6t
Xbit_r94_c252 bl_252 br_252 wl_94 vdd gnd cell_6t
Xbit_r95_c252 bl_252 br_252 wl_95 vdd gnd cell_6t
Xbit_r96_c252 bl_252 br_252 wl_96 vdd gnd cell_6t
Xbit_r97_c252 bl_252 br_252 wl_97 vdd gnd cell_6t
Xbit_r98_c252 bl_252 br_252 wl_98 vdd gnd cell_6t
Xbit_r99_c252 bl_252 br_252 wl_99 vdd gnd cell_6t
Xbit_r100_c252 bl_252 br_252 wl_100 vdd gnd cell_6t
Xbit_r101_c252 bl_252 br_252 wl_101 vdd gnd cell_6t
Xbit_r102_c252 bl_252 br_252 wl_102 vdd gnd cell_6t
Xbit_r103_c252 bl_252 br_252 wl_103 vdd gnd cell_6t
Xbit_r104_c252 bl_252 br_252 wl_104 vdd gnd cell_6t
Xbit_r105_c252 bl_252 br_252 wl_105 vdd gnd cell_6t
Xbit_r106_c252 bl_252 br_252 wl_106 vdd gnd cell_6t
Xbit_r107_c252 bl_252 br_252 wl_107 vdd gnd cell_6t
Xbit_r108_c252 bl_252 br_252 wl_108 vdd gnd cell_6t
Xbit_r109_c252 bl_252 br_252 wl_109 vdd gnd cell_6t
Xbit_r110_c252 bl_252 br_252 wl_110 vdd gnd cell_6t
Xbit_r111_c252 bl_252 br_252 wl_111 vdd gnd cell_6t
Xbit_r112_c252 bl_252 br_252 wl_112 vdd gnd cell_6t
Xbit_r113_c252 bl_252 br_252 wl_113 vdd gnd cell_6t
Xbit_r114_c252 bl_252 br_252 wl_114 vdd gnd cell_6t
Xbit_r115_c252 bl_252 br_252 wl_115 vdd gnd cell_6t
Xbit_r116_c252 bl_252 br_252 wl_116 vdd gnd cell_6t
Xbit_r117_c252 bl_252 br_252 wl_117 vdd gnd cell_6t
Xbit_r118_c252 bl_252 br_252 wl_118 vdd gnd cell_6t
Xbit_r119_c252 bl_252 br_252 wl_119 vdd gnd cell_6t
Xbit_r120_c252 bl_252 br_252 wl_120 vdd gnd cell_6t
Xbit_r121_c252 bl_252 br_252 wl_121 vdd gnd cell_6t
Xbit_r122_c252 bl_252 br_252 wl_122 vdd gnd cell_6t
Xbit_r123_c252 bl_252 br_252 wl_123 vdd gnd cell_6t
Xbit_r124_c252 bl_252 br_252 wl_124 vdd gnd cell_6t
Xbit_r125_c252 bl_252 br_252 wl_125 vdd gnd cell_6t
Xbit_r126_c252 bl_252 br_252 wl_126 vdd gnd cell_6t
Xbit_r127_c252 bl_252 br_252 wl_127 vdd gnd cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd cell_6t
Xbit_r1_c253 bl_253 br_253 wl_1 vdd gnd cell_6t
Xbit_r2_c253 bl_253 br_253 wl_2 vdd gnd cell_6t
Xbit_r3_c253 bl_253 br_253 wl_3 vdd gnd cell_6t
Xbit_r4_c253 bl_253 br_253 wl_4 vdd gnd cell_6t
Xbit_r5_c253 bl_253 br_253 wl_5 vdd gnd cell_6t
Xbit_r6_c253 bl_253 br_253 wl_6 vdd gnd cell_6t
Xbit_r7_c253 bl_253 br_253 wl_7 vdd gnd cell_6t
Xbit_r8_c253 bl_253 br_253 wl_8 vdd gnd cell_6t
Xbit_r9_c253 bl_253 br_253 wl_9 vdd gnd cell_6t
Xbit_r10_c253 bl_253 br_253 wl_10 vdd gnd cell_6t
Xbit_r11_c253 bl_253 br_253 wl_11 vdd gnd cell_6t
Xbit_r12_c253 bl_253 br_253 wl_12 vdd gnd cell_6t
Xbit_r13_c253 bl_253 br_253 wl_13 vdd gnd cell_6t
Xbit_r14_c253 bl_253 br_253 wl_14 vdd gnd cell_6t
Xbit_r15_c253 bl_253 br_253 wl_15 vdd gnd cell_6t
Xbit_r16_c253 bl_253 br_253 wl_16 vdd gnd cell_6t
Xbit_r17_c253 bl_253 br_253 wl_17 vdd gnd cell_6t
Xbit_r18_c253 bl_253 br_253 wl_18 vdd gnd cell_6t
Xbit_r19_c253 bl_253 br_253 wl_19 vdd gnd cell_6t
Xbit_r20_c253 bl_253 br_253 wl_20 vdd gnd cell_6t
Xbit_r21_c253 bl_253 br_253 wl_21 vdd gnd cell_6t
Xbit_r22_c253 bl_253 br_253 wl_22 vdd gnd cell_6t
Xbit_r23_c253 bl_253 br_253 wl_23 vdd gnd cell_6t
Xbit_r24_c253 bl_253 br_253 wl_24 vdd gnd cell_6t
Xbit_r25_c253 bl_253 br_253 wl_25 vdd gnd cell_6t
Xbit_r26_c253 bl_253 br_253 wl_26 vdd gnd cell_6t
Xbit_r27_c253 bl_253 br_253 wl_27 vdd gnd cell_6t
Xbit_r28_c253 bl_253 br_253 wl_28 vdd gnd cell_6t
Xbit_r29_c253 bl_253 br_253 wl_29 vdd gnd cell_6t
Xbit_r30_c253 bl_253 br_253 wl_30 vdd gnd cell_6t
Xbit_r31_c253 bl_253 br_253 wl_31 vdd gnd cell_6t
Xbit_r32_c253 bl_253 br_253 wl_32 vdd gnd cell_6t
Xbit_r33_c253 bl_253 br_253 wl_33 vdd gnd cell_6t
Xbit_r34_c253 bl_253 br_253 wl_34 vdd gnd cell_6t
Xbit_r35_c253 bl_253 br_253 wl_35 vdd gnd cell_6t
Xbit_r36_c253 bl_253 br_253 wl_36 vdd gnd cell_6t
Xbit_r37_c253 bl_253 br_253 wl_37 vdd gnd cell_6t
Xbit_r38_c253 bl_253 br_253 wl_38 vdd gnd cell_6t
Xbit_r39_c253 bl_253 br_253 wl_39 vdd gnd cell_6t
Xbit_r40_c253 bl_253 br_253 wl_40 vdd gnd cell_6t
Xbit_r41_c253 bl_253 br_253 wl_41 vdd gnd cell_6t
Xbit_r42_c253 bl_253 br_253 wl_42 vdd gnd cell_6t
Xbit_r43_c253 bl_253 br_253 wl_43 vdd gnd cell_6t
Xbit_r44_c253 bl_253 br_253 wl_44 vdd gnd cell_6t
Xbit_r45_c253 bl_253 br_253 wl_45 vdd gnd cell_6t
Xbit_r46_c253 bl_253 br_253 wl_46 vdd gnd cell_6t
Xbit_r47_c253 bl_253 br_253 wl_47 vdd gnd cell_6t
Xbit_r48_c253 bl_253 br_253 wl_48 vdd gnd cell_6t
Xbit_r49_c253 bl_253 br_253 wl_49 vdd gnd cell_6t
Xbit_r50_c253 bl_253 br_253 wl_50 vdd gnd cell_6t
Xbit_r51_c253 bl_253 br_253 wl_51 vdd gnd cell_6t
Xbit_r52_c253 bl_253 br_253 wl_52 vdd gnd cell_6t
Xbit_r53_c253 bl_253 br_253 wl_53 vdd gnd cell_6t
Xbit_r54_c253 bl_253 br_253 wl_54 vdd gnd cell_6t
Xbit_r55_c253 bl_253 br_253 wl_55 vdd gnd cell_6t
Xbit_r56_c253 bl_253 br_253 wl_56 vdd gnd cell_6t
Xbit_r57_c253 bl_253 br_253 wl_57 vdd gnd cell_6t
Xbit_r58_c253 bl_253 br_253 wl_58 vdd gnd cell_6t
Xbit_r59_c253 bl_253 br_253 wl_59 vdd gnd cell_6t
Xbit_r60_c253 bl_253 br_253 wl_60 vdd gnd cell_6t
Xbit_r61_c253 bl_253 br_253 wl_61 vdd gnd cell_6t
Xbit_r62_c253 bl_253 br_253 wl_62 vdd gnd cell_6t
Xbit_r63_c253 bl_253 br_253 wl_63 vdd gnd cell_6t
Xbit_r64_c253 bl_253 br_253 wl_64 vdd gnd cell_6t
Xbit_r65_c253 bl_253 br_253 wl_65 vdd gnd cell_6t
Xbit_r66_c253 bl_253 br_253 wl_66 vdd gnd cell_6t
Xbit_r67_c253 bl_253 br_253 wl_67 vdd gnd cell_6t
Xbit_r68_c253 bl_253 br_253 wl_68 vdd gnd cell_6t
Xbit_r69_c253 bl_253 br_253 wl_69 vdd gnd cell_6t
Xbit_r70_c253 bl_253 br_253 wl_70 vdd gnd cell_6t
Xbit_r71_c253 bl_253 br_253 wl_71 vdd gnd cell_6t
Xbit_r72_c253 bl_253 br_253 wl_72 vdd gnd cell_6t
Xbit_r73_c253 bl_253 br_253 wl_73 vdd gnd cell_6t
Xbit_r74_c253 bl_253 br_253 wl_74 vdd gnd cell_6t
Xbit_r75_c253 bl_253 br_253 wl_75 vdd gnd cell_6t
Xbit_r76_c253 bl_253 br_253 wl_76 vdd gnd cell_6t
Xbit_r77_c253 bl_253 br_253 wl_77 vdd gnd cell_6t
Xbit_r78_c253 bl_253 br_253 wl_78 vdd gnd cell_6t
Xbit_r79_c253 bl_253 br_253 wl_79 vdd gnd cell_6t
Xbit_r80_c253 bl_253 br_253 wl_80 vdd gnd cell_6t
Xbit_r81_c253 bl_253 br_253 wl_81 vdd gnd cell_6t
Xbit_r82_c253 bl_253 br_253 wl_82 vdd gnd cell_6t
Xbit_r83_c253 bl_253 br_253 wl_83 vdd gnd cell_6t
Xbit_r84_c253 bl_253 br_253 wl_84 vdd gnd cell_6t
Xbit_r85_c253 bl_253 br_253 wl_85 vdd gnd cell_6t
Xbit_r86_c253 bl_253 br_253 wl_86 vdd gnd cell_6t
Xbit_r87_c253 bl_253 br_253 wl_87 vdd gnd cell_6t
Xbit_r88_c253 bl_253 br_253 wl_88 vdd gnd cell_6t
Xbit_r89_c253 bl_253 br_253 wl_89 vdd gnd cell_6t
Xbit_r90_c253 bl_253 br_253 wl_90 vdd gnd cell_6t
Xbit_r91_c253 bl_253 br_253 wl_91 vdd gnd cell_6t
Xbit_r92_c253 bl_253 br_253 wl_92 vdd gnd cell_6t
Xbit_r93_c253 bl_253 br_253 wl_93 vdd gnd cell_6t
Xbit_r94_c253 bl_253 br_253 wl_94 vdd gnd cell_6t
Xbit_r95_c253 bl_253 br_253 wl_95 vdd gnd cell_6t
Xbit_r96_c253 bl_253 br_253 wl_96 vdd gnd cell_6t
Xbit_r97_c253 bl_253 br_253 wl_97 vdd gnd cell_6t
Xbit_r98_c253 bl_253 br_253 wl_98 vdd gnd cell_6t
Xbit_r99_c253 bl_253 br_253 wl_99 vdd gnd cell_6t
Xbit_r100_c253 bl_253 br_253 wl_100 vdd gnd cell_6t
Xbit_r101_c253 bl_253 br_253 wl_101 vdd gnd cell_6t
Xbit_r102_c253 bl_253 br_253 wl_102 vdd gnd cell_6t
Xbit_r103_c253 bl_253 br_253 wl_103 vdd gnd cell_6t
Xbit_r104_c253 bl_253 br_253 wl_104 vdd gnd cell_6t
Xbit_r105_c253 bl_253 br_253 wl_105 vdd gnd cell_6t
Xbit_r106_c253 bl_253 br_253 wl_106 vdd gnd cell_6t
Xbit_r107_c253 bl_253 br_253 wl_107 vdd gnd cell_6t
Xbit_r108_c253 bl_253 br_253 wl_108 vdd gnd cell_6t
Xbit_r109_c253 bl_253 br_253 wl_109 vdd gnd cell_6t
Xbit_r110_c253 bl_253 br_253 wl_110 vdd gnd cell_6t
Xbit_r111_c253 bl_253 br_253 wl_111 vdd gnd cell_6t
Xbit_r112_c253 bl_253 br_253 wl_112 vdd gnd cell_6t
Xbit_r113_c253 bl_253 br_253 wl_113 vdd gnd cell_6t
Xbit_r114_c253 bl_253 br_253 wl_114 vdd gnd cell_6t
Xbit_r115_c253 bl_253 br_253 wl_115 vdd gnd cell_6t
Xbit_r116_c253 bl_253 br_253 wl_116 vdd gnd cell_6t
Xbit_r117_c253 bl_253 br_253 wl_117 vdd gnd cell_6t
Xbit_r118_c253 bl_253 br_253 wl_118 vdd gnd cell_6t
Xbit_r119_c253 bl_253 br_253 wl_119 vdd gnd cell_6t
Xbit_r120_c253 bl_253 br_253 wl_120 vdd gnd cell_6t
Xbit_r121_c253 bl_253 br_253 wl_121 vdd gnd cell_6t
Xbit_r122_c253 bl_253 br_253 wl_122 vdd gnd cell_6t
Xbit_r123_c253 bl_253 br_253 wl_123 vdd gnd cell_6t
Xbit_r124_c253 bl_253 br_253 wl_124 vdd gnd cell_6t
Xbit_r125_c253 bl_253 br_253 wl_125 vdd gnd cell_6t
Xbit_r126_c253 bl_253 br_253 wl_126 vdd gnd cell_6t
Xbit_r127_c253 bl_253 br_253 wl_127 vdd gnd cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd cell_6t
Xbit_r1_c254 bl_254 br_254 wl_1 vdd gnd cell_6t
Xbit_r2_c254 bl_254 br_254 wl_2 vdd gnd cell_6t
Xbit_r3_c254 bl_254 br_254 wl_3 vdd gnd cell_6t
Xbit_r4_c254 bl_254 br_254 wl_4 vdd gnd cell_6t
Xbit_r5_c254 bl_254 br_254 wl_5 vdd gnd cell_6t
Xbit_r6_c254 bl_254 br_254 wl_6 vdd gnd cell_6t
Xbit_r7_c254 bl_254 br_254 wl_7 vdd gnd cell_6t
Xbit_r8_c254 bl_254 br_254 wl_8 vdd gnd cell_6t
Xbit_r9_c254 bl_254 br_254 wl_9 vdd gnd cell_6t
Xbit_r10_c254 bl_254 br_254 wl_10 vdd gnd cell_6t
Xbit_r11_c254 bl_254 br_254 wl_11 vdd gnd cell_6t
Xbit_r12_c254 bl_254 br_254 wl_12 vdd gnd cell_6t
Xbit_r13_c254 bl_254 br_254 wl_13 vdd gnd cell_6t
Xbit_r14_c254 bl_254 br_254 wl_14 vdd gnd cell_6t
Xbit_r15_c254 bl_254 br_254 wl_15 vdd gnd cell_6t
Xbit_r16_c254 bl_254 br_254 wl_16 vdd gnd cell_6t
Xbit_r17_c254 bl_254 br_254 wl_17 vdd gnd cell_6t
Xbit_r18_c254 bl_254 br_254 wl_18 vdd gnd cell_6t
Xbit_r19_c254 bl_254 br_254 wl_19 vdd gnd cell_6t
Xbit_r20_c254 bl_254 br_254 wl_20 vdd gnd cell_6t
Xbit_r21_c254 bl_254 br_254 wl_21 vdd gnd cell_6t
Xbit_r22_c254 bl_254 br_254 wl_22 vdd gnd cell_6t
Xbit_r23_c254 bl_254 br_254 wl_23 vdd gnd cell_6t
Xbit_r24_c254 bl_254 br_254 wl_24 vdd gnd cell_6t
Xbit_r25_c254 bl_254 br_254 wl_25 vdd gnd cell_6t
Xbit_r26_c254 bl_254 br_254 wl_26 vdd gnd cell_6t
Xbit_r27_c254 bl_254 br_254 wl_27 vdd gnd cell_6t
Xbit_r28_c254 bl_254 br_254 wl_28 vdd gnd cell_6t
Xbit_r29_c254 bl_254 br_254 wl_29 vdd gnd cell_6t
Xbit_r30_c254 bl_254 br_254 wl_30 vdd gnd cell_6t
Xbit_r31_c254 bl_254 br_254 wl_31 vdd gnd cell_6t
Xbit_r32_c254 bl_254 br_254 wl_32 vdd gnd cell_6t
Xbit_r33_c254 bl_254 br_254 wl_33 vdd gnd cell_6t
Xbit_r34_c254 bl_254 br_254 wl_34 vdd gnd cell_6t
Xbit_r35_c254 bl_254 br_254 wl_35 vdd gnd cell_6t
Xbit_r36_c254 bl_254 br_254 wl_36 vdd gnd cell_6t
Xbit_r37_c254 bl_254 br_254 wl_37 vdd gnd cell_6t
Xbit_r38_c254 bl_254 br_254 wl_38 vdd gnd cell_6t
Xbit_r39_c254 bl_254 br_254 wl_39 vdd gnd cell_6t
Xbit_r40_c254 bl_254 br_254 wl_40 vdd gnd cell_6t
Xbit_r41_c254 bl_254 br_254 wl_41 vdd gnd cell_6t
Xbit_r42_c254 bl_254 br_254 wl_42 vdd gnd cell_6t
Xbit_r43_c254 bl_254 br_254 wl_43 vdd gnd cell_6t
Xbit_r44_c254 bl_254 br_254 wl_44 vdd gnd cell_6t
Xbit_r45_c254 bl_254 br_254 wl_45 vdd gnd cell_6t
Xbit_r46_c254 bl_254 br_254 wl_46 vdd gnd cell_6t
Xbit_r47_c254 bl_254 br_254 wl_47 vdd gnd cell_6t
Xbit_r48_c254 bl_254 br_254 wl_48 vdd gnd cell_6t
Xbit_r49_c254 bl_254 br_254 wl_49 vdd gnd cell_6t
Xbit_r50_c254 bl_254 br_254 wl_50 vdd gnd cell_6t
Xbit_r51_c254 bl_254 br_254 wl_51 vdd gnd cell_6t
Xbit_r52_c254 bl_254 br_254 wl_52 vdd gnd cell_6t
Xbit_r53_c254 bl_254 br_254 wl_53 vdd gnd cell_6t
Xbit_r54_c254 bl_254 br_254 wl_54 vdd gnd cell_6t
Xbit_r55_c254 bl_254 br_254 wl_55 vdd gnd cell_6t
Xbit_r56_c254 bl_254 br_254 wl_56 vdd gnd cell_6t
Xbit_r57_c254 bl_254 br_254 wl_57 vdd gnd cell_6t
Xbit_r58_c254 bl_254 br_254 wl_58 vdd gnd cell_6t
Xbit_r59_c254 bl_254 br_254 wl_59 vdd gnd cell_6t
Xbit_r60_c254 bl_254 br_254 wl_60 vdd gnd cell_6t
Xbit_r61_c254 bl_254 br_254 wl_61 vdd gnd cell_6t
Xbit_r62_c254 bl_254 br_254 wl_62 vdd gnd cell_6t
Xbit_r63_c254 bl_254 br_254 wl_63 vdd gnd cell_6t
Xbit_r64_c254 bl_254 br_254 wl_64 vdd gnd cell_6t
Xbit_r65_c254 bl_254 br_254 wl_65 vdd gnd cell_6t
Xbit_r66_c254 bl_254 br_254 wl_66 vdd gnd cell_6t
Xbit_r67_c254 bl_254 br_254 wl_67 vdd gnd cell_6t
Xbit_r68_c254 bl_254 br_254 wl_68 vdd gnd cell_6t
Xbit_r69_c254 bl_254 br_254 wl_69 vdd gnd cell_6t
Xbit_r70_c254 bl_254 br_254 wl_70 vdd gnd cell_6t
Xbit_r71_c254 bl_254 br_254 wl_71 vdd gnd cell_6t
Xbit_r72_c254 bl_254 br_254 wl_72 vdd gnd cell_6t
Xbit_r73_c254 bl_254 br_254 wl_73 vdd gnd cell_6t
Xbit_r74_c254 bl_254 br_254 wl_74 vdd gnd cell_6t
Xbit_r75_c254 bl_254 br_254 wl_75 vdd gnd cell_6t
Xbit_r76_c254 bl_254 br_254 wl_76 vdd gnd cell_6t
Xbit_r77_c254 bl_254 br_254 wl_77 vdd gnd cell_6t
Xbit_r78_c254 bl_254 br_254 wl_78 vdd gnd cell_6t
Xbit_r79_c254 bl_254 br_254 wl_79 vdd gnd cell_6t
Xbit_r80_c254 bl_254 br_254 wl_80 vdd gnd cell_6t
Xbit_r81_c254 bl_254 br_254 wl_81 vdd gnd cell_6t
Xbit_r82_c254 bl_254 br_254 wl_82 vdd gnd cell_6t
Xbit_r83_c254 bl_254 br_254 wl_83 vdd gnd cell_6t
Xbit_r84_c254 bl_254 br_254 wl_84 vdd gnd cell_6t
Xbit_r85_c254 bl_254 br_254 wl_85 vdd gnd cell_6t
Xbit_r86_c254 bl_254 br_254 wl_86 vdd gnd cell_6t
Xbit_r87_c254 bl_254 br_254 wl_87 vdd gnd cell_6t
Xbit_r88_c254 bl_254 br_254 wl_88 vdd gnd cell_6t
Xbit_r89_c254 bl_254 br_254 wl_89 vdd gnd cell_6t
Xbit_r90_c254 bl_254 br_254 wl_90 vdd gnd cell_6t
Xbit_r91_c254 bl_254 br_254 wl_91 vdd gnd cell_6t
Xbit_r92_c254 bl_254 br_254 wl_92 vdd gnd cell_6t
Xbit_r93_c254 bl_254 br_254 wl_93 vdd gnd cell_6t
Xbit_r94_c254 bl_254 br_254 wl_94 vdd gnd cell_6t
Xbit_r95_c254 bl_254 br_254 wl_95 vdd gnd cell_6t
Xbit_r96_c254 bl_254 br_254 wl_96 vdd gnd cell_6t
Xbit_r97_c254 bl_254 br_254 wl_97 vdd gnd cell_6t
Xbit_r98_c254 bl_254 br_254 wl_98 vdd gnd cell_6t
Xbit_r99_c254 bl_254 br_254 wl_99 vdd gnd cell_6t
Xbit_r100_c254 bl_254 br_254 wl_100 vdd gnd cell_6t
Xbit_r101_c254 bl_254 br_254 wl_101 vdd gnd cell_6t
Xbit_r102_c254 bl_254 br_254 wl_102 vdd gnd cell_6t
Xbit_r103_c254 bl_254 br_254 wl_103 vdd gnd cell_6t
Xbit_r104_c254 bl_254 br_254 wl_104 vdd gnd cell_6t
Xbit_r105_c254 bl_254 br_254 wl_105 vdd gnd cell_6t
Xbit_r106_c254 bl_254 br_254 wl_106 vdd gnd cell_6t
Xbit_r107_c254 bl_254 br_254 wl_107 vdd gnd cell_6t
Xbit_r108_c254 bl_254 br_254 wl_108 vdd gnd cell_6t
Xbit_r109_c254 bl_254 br_254 wl_109 vdd gnd cell_6t
Xbit_r110_c254 bl_254 br_254 wl_110 vdd gnd cell_6t
Xbit_r111_c254 bl_254 br_254 wl_111 vdd gnd cell_6t
Xbit_r112_c254 bl_254 br_254 wl_112 vdd gnd cell_6t
Xbit_r113_c254 bl_254 br_254 wl_113 vdd gnd cell_6t
Xbit_r114_c254 bl_254 br_254 wl_114 vdd gnd cell_6t
Xbit_r115_c254 bl_254 br_254 wl_115 vdd gnd cell_6t
Xbit_r116_c254 bl_254 br_254 wl_116 vdd gnd cell_6t
Xbit_r117_c254 bl_254 br_254 wl_117 vdd gnd cell_6t
Xbit_r118_c254 bl_254 br_254 wl_118 vdd gnd cell_6t
Xbit_r119_c254 bl_254 br_254 wl_119 vdd gnd cell_6t
Xbit_r120_c254 bl_254 br_254 wl_120 vdd gnd cell_6t
Xbit_r121_c254 bl_254 br_254 wl_121 vdd gnd cell_6t
Xbit_r122_c254 bl_254 br_254 wl_122 vdd gnd cell_6t
Xbit_r123_c254 bl_254 br_254 wl_123 vdd gnd cell_6t
Xbit_r124_c254 bl_254 br_254 wl_124 vdd gnd cell_6t
Xbit_r125_c254 bl_254 br_254 wl_125 vdd gnd cell_6t
Xbit_r126_c254 bl_254 br_254 wl_126 vdd gnd cell_6t
Xbit_r127_c254 bl_254 br_254 wl_127 vdd gnd cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd cell_6t
Xbit_r1_c255 bl_255 br_255 wl_1 vdd gnd cell_6t
Xbit_r2_c255 bl_255 br_255 wl_2 vdd gnd cell_6t
Xbit_r3_c255 bl_255 br_255 wl_3 vdd gnd cell_6t
Xbit_r4_c255 bl_255 br_255 wl_4 vdd gnd cell_6t
Xbit_r5_c255 bl_255 br_255 wl_5 vdd gnd cell_6t
Xbit_r6_c255 bl_255 br_255 wl_6 vdd gnd cell_6t
Xbit_r7_c255 bl_255 br_255 wl_7 vdd gnd cell_6t
Xbit_r8_c255 bl_255 br_255 wl_8 vdd gnd cell_6t
Xbit_r9_c255 bl_255 br_255 wl_9 vdd gnd cell_6t
Xbit_r10_c255 bl_255 br_255 wl_10 vdd gnd cell_6t
Xbit_r11_c255 bl_255 br_255 wl_11 vdd gnd cell_6t
Xbit_r12_c255 bl_255 br_255 wl_12 vdd gnd cell_6t
Xbit_r13_c255 bl_255 br_255 wl_13 vdd gnd cell_6t
Xbit_r14_c255 bl_255 br_255 wl_14 vdd gnd cell_6t
Xbit_r15_c255 bl_255 br_255 wl_15 vdd gnd cell_6t
Xbit_r16_c255 bl_255 br_255 wl_16 vdd gnd cell_6t
Xbit_r17_c255 bl_255 br_255 wl_17 vdd gnd cell_6t
Xbit_r18_c255 bl_255 br_255 wl_18 vdd gnd cell_6t
Xbit_r19_c255 bl_255 br_255 wl_19 vdd gnd cell_6t
Xbit_r20_c255 bl_255 br_255 wl_20 vdd gnd cell_6t
Xbit_r21_c255 bl_255 br_255 wl_21 vdd gnd cell_6t
Xbit_r22_c255 bl_255 br_255 wl_22 vdd gnd cell_6t
Xbit_r23_c255 bl_255 br_255 wl_23 vdd gnd cell_6t
Xbit_r24_c255 bl_255 br_255 wl_24 vdd gnd cell_6t
Xbit_r25_c255 bl_255 br_255 wl_25 vdd gnd cell_6t
Xbit_r26_c255 bl_255 br_255 wl_26 vdd gnd cell_6t
Xbit_r27_c255 bl_255 br_255 wl_27 vdd gnd cell_6t
Xbit_r28_c255 bl_255 br_255 wl_28 vdd gnd cell_6t
Xbit_r29_c255 bl_255 br_255 wl_29 vdd gnd cell_6t
Xbit_r30_c255 bl_255 br_255 wl_30 vdd gnd cell_6t
Xbit_r31_c255 bl_255 br_255 wl_31 vdd gnd cell_6t
Xbit_r32_c255 bl_255 br_255 wl_32 vdd gnd cell_6t
Xbit_r33_c255 bl_255 br_255 wl_33 vdd gnd cell_6t
Xbit_r34_c255 bl_255 br_255 wl_34 vdd gnd cell_6t
Xbit_r35_c255 bl_255 br_255 wl_35 vdd gnd cell_6t
Xbit_r36_c255 bl_255 br_255 wl_36 vdd gnd cell_6t
Xbit_r37_c255 bl_255 br_255 wl_37 vdd gnd cell_6t
Xbit_r38_c255 bl_255 br_255 wl_38 vdd gnd cell_6t
Xbit_r39_c255 bl_255 br_255 wl_39 vdd gnd cell_6t
Xbit_r40_c255 bl_255 br_255 wl_40 vdd gnd cell_6t
Xbit_r41_c255 bl_255 br_255 wl_41 vdd gnd cell_6t
Xbit_r42_c255 bl_255 br_255 wl_42 vdd gnd cell_6t
Xbit_r43_c255 bl_255 br_255 wl_43 vdd gnd cell_6t
Xbit_r44_c255 bl_255 br_255 wl_44 vdd gnd cell_6t
Xbit_r45_c255 bl_255 br_255 wl_45 vdd gnd cell_6t
Xbit_r46_c255 bl_255 br_255 wl_46 vdd gnd cell_6t
Xbit_r47_c255 bl_255 br_255 wl_47 vdd gnd cell_6t
Xbit_r48_c255 bl_255 br_255 wl_48 vdd gnd cell_6t
Xbit_r49_c255 bl_255 br_255 wl_49 vdd gnd cell_6t
Xbit_r50_c255 bl_255 br_255 wl_50 vdd gnd cell_6t
Xbit_r51_c255 bl_255 br_255 wl_51 vdd gnd cell_6t
Xbit_r52_c255 bl_255 br_255 wl_52 vdd gnd cell_6t
Xbit_r53_c255 bl_255 br_255 wl_53 vdd gnd cell_6t
Xbit_r54_c255 bl_255 br_255 wl_54 vdd gnd cell_6t
Xbit_r55_c255 bl_255 br_255 wl_55 vdd gnd cell_6t
Xbit_r56_c255 bl_255 br_255 wl_56 vdd gnd cell_6t
Xbit_r57_c255 bl_255 br_255 wl_57 vdd gnd cell_6t
Xbit_r58_c255 bl_255 br_255 wl_58 vdd gnd cell_6t
Xbit_r59_c255 bl_255 br_255 wl_59 vdd gnd cell_6t
Xbit_r60_c255 bl_255 br_255 wl_60 vdd gnd cell_6t
Xbit_r61_c255 bl_255 br_255 wl_61 vdd gnd cell_6t
Xbit_r62_c255 bl_255 br_255 wl_62 vdd gnd cell_6t
Xbit_r63_c255 bl_255 br_255 wl_63 vdd gnd cell_6t
Xbit_r64_c255 bl_255 br_255 wl_64 vdd gnd cell_6t
Xbit_r65_c255 bl_255 br_255 wl_65 vdd gnd cell_6t
Xbit_r66_c255 bl_255 br_255 wl_66 vdd gnd cell_6t
Xbit_r67_c255 bl_255 br_255 wl_67 vdd gnd cell_6t
Xbit_r68_c255 bl_255 br_255 wl_68 vdd gnd cell_6t
Xbit_r69_c255 bl_255 br_255 wl_69 vdd gnd cell_6t
Xbit_r70_c255 bl_255 br_255 wl_70 vdd gnd cell_6t
Xbit_r71_c255 bl_255 br_255 wl_71 vdd gnd cell_6t
Xbit_r72_c255 bl_255 br_255 wl_72 vdd gnd cell_6t
Xbit_r73_c255 bl_255 br_255 wl_73 vdd gnd cell_6t
Xbit_r74_c255 bl_255 br_255 wl_74 vdd gnd cell_6t
Xbit_r75_c255 bl_255 br_255 wl_75 vdd gnd cell_6t
Xbit_r76_c255 bl_255 br_255 wl_76 vdd gnd cell_6t
Xbit_r77_c255 bl_255 br_255 wl_77 vdd gnd cell_6t
Xbit_r78_c255 bl_255 br_255 wl_78 vdd gnd cell_6t
Xbit_r79_c255 bl_255 br_255 wl_79 vdd gnd cell_6t
Xbit_r80_c255 bl_255 br_255 wl_80 vdd gnd cell_6t
Xbit_r81_c255 bl_255 br_255 wl_81 vdd gnd cell_6t
Xbit_r82_c255 bl_255 br_255 wl_82 vdd gnd cell_6t
Xbit_r83_c255 bl_255 br_255 wl_83 vdd gnd cell_6t
Xbit_r84_c255 bl_255 br_255 wl_84 vdd gnd cell_6t
Xbit_r85_c255 bl_255 br_255 wl_85 vdd gnd cell_6t
Xbit_r86_c255 bl_255 br_255 wl_86 vdd gnd cell_6t
Xbit_r87_c255 bl_255 br_255 wl_87 vdd gnd cell_6t
Xbit_r88_c255 bl_255 br_255 wl_88 vdd gnd cell_6t
Xbit_r89_c255 bl_255 br_255 wl_89 vdd gnd cell_6t
Xbit_r90_c255 bl_255 br_255 wl_90 vdd gnd cell_6t
Xbit_r91_c255 bl_255 br_255 wl_91 vdd gnd cell_6t
Xbit_r92_c255 bl_255 br_255 wl_92 vdd gnd cell_6t
Xbit_r93_c255 bl_255 br_255 wl_93 vdd gnd cell_6t
Xbit_r94_c255 bl_255 br_255 wl_94 vdd gnd cell_6t
Xbit_r95_c255 bl_255 br_255 wl_95 vdd gnd cell_6t
Xbit_r96_c255 bl_255 br_255 wl_96 vdd gnd cell_6t
Xbit_r97_c255 bl_255 br_255 wl_97 vdd gnd cell_6t
Xbit_r98_c255 bl_255 br_255 wl_98 vdd gnd cell_6t
Xbit_r99_c255 bl_255 br_255 wl_99 vdd gnd cell_6t
Xbit_r100_c255 bl_255 br_255 wl_100 vdd gnd cell_6t
Xbit_r101_c255 bl_255 br_255 wl_101 vdd gnd cell_6t
Xbit_r102_c255 bl_255 br_255 wl_102 vdd gnd cell_6t
Xbit_r103_c255 bl_255 br_255 wl_103 vdd gnd cell_6t
Xbit_r104_c255 bl_255 br_255 wl_104 vdd gnd cell_6t
Xbit_r105_c255 bl_255 br_255 wl_105 vdd gnd cell_6t
Xbit_r106_c255 bl_255 br_255 wl_106 vdd gnd cell_6t
Xbit_r107_c255 bl_255 br_255 wl_107 vdd gnd cell_6t
Xbit_r108_c255 bl_255 br_255 wl_108 vdd gnd cell_6t
Xbit_r109_c255 bl_255 br_255 wl_109 vdd gnd cell_6t
Xbit_r110_c255 bl_255 br_255 wl_110 vdd gnd cell_6t
Xbit_r111_c255 bl_255 br_255 wl_111 vdd gnd cell_6t
Xbit_r112_c255 bl_255 br_255 wl_112 vdd gnd cell_6t
Xbit_r113_c255 bl_255 br_255 wl_113 vdd gnd cell_6t
Xbit_r114_c255 bl_255 br_255 wl_114 vdd gnd cell_6t
Xbit_r115_c255 bl_255 br_255 wl_115 vdd gnd cell_6t
Xbit_r116_c255 bl_255 br_255 wl_116 vdd gnd cell_6t
Xbit_r117_c255 bl_255 br_255 wl_117 vdd gnd cell_6t
Xbit_r118_c255 bl_255 br_255 wl_118 vdd gnd cell_6t
Xbit_r119_c255 bl_255 br_255 wl_119 vdd gnd cell_6t
Xbit_r120_c255 bl_255 br_255 wl_120 vdd gnd cell_6t
Xbit_r121_c255 bl_255 br_255 wl_121 vdd gnd cell_6t
Xbit_r122_c255 bl_255 br_255 wl_122 vdd gnd cell_6t
Xbit_r123_c255 bl_255 br_255 wl_123 vdd gnd cell_6t
Xbit_r124_c255 bl_255 br_255 wl_124 vdd gnd cell_6t
Xbit_r125_c255 bl_255 br_255 wl_125 vdd gnd cell_6t
Xbit_r126_c255 bl_255 br_255 wl_126 vdd gnd cell_6t
Xbit_r127_c255 bl_255 br_255 wl_127 vdd gnd cell_6t
.ENDS bitcell_array_0

.SUBCKT replica_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 vdd Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 vdd Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q vdd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q vdd vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br wl vdd gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT dummy_cell_6t bl br wl vdd gnd
* Inverter 1
MM0 Qbar Q gnd gnd NMOS_VTG W=205.00n L=50n
MM4 Qbar Q vdd vdd PMOS_VTG W=90n L=50n

* Inverer 2
MM1 Q Qbar gnd gnd NMOS_VTG W=205.00n L=50n
MM5 Q Qbar vdd vdd PMOS_VTG W=90n L=50n

* Access transistors
MM3 bl_noconn wl Q gnd NMOS_VTG W=135.00n L=50n
MM2 br_noconn wl Qbar gnd NMOS_VTG W=135.00n L=50n
.ENDS cell_6t


.SUBCKT replica_column_0 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 vdd gnd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xrbc_1 bl_0 br_0 wl_1 vdd gnd replica_cell_6t
Xrbc_2 bl_0 br_0 wl_2 vdd gnd replica_cell_6t
Xrbc_3 bl_0 br_0 wl_3 vdd gnd replica_cell_6t
Xrbc_4 bl_0 br_0 wl_4 vdd gnd replica_cell_6t
Xrbc_5 bl_0 br_0 wl_5 vdd gnd replica_cell_6t
Xrbc_6 bl_0 br_0 wl_6 vdd gnd replica_cell_6t
Xrbc_7 bl_0 br_0 wl_7 vdd gnd replica_cell_6t
Xrbc_8 bl_0 br_0 wl_8 vdd gnd replica_cell_6t
Xrbc_9 bl_0 br_0 wl_9 vdd gnd replica_cell_6t
Xrbc_10 bl_0 br_0 wl_10 vdd gnd replica_cell_6t
Xrbc_11 bl_0 br_0 wl_11 vdd gnd replica_cell_6t
Xrbc_12 bl_0 br_0 wl_12 vdd gnd replica_cell_6t
Xrbc_13 bl_0 br_0 wl_13 vdd gnd replica_cell_6t
Xrbc_14 bl_0 br_0 wl_14 vdd gnd replica_cell_6t
Xrbc_15 bl_0 br_0 wl_15 vdd gnd replica_cell_6t
Xrbc_16 bl_0 br_0 wl_16 vdd gnd replica_cell_6t
Xrbc_17 bl_0 br_0 wl_17 vdd gnd replica_cell_6t
Xrbc_18 bl_0 br_0 wl_18 vdd gnd replica_cell_6t
Xrbc_19 bl_0 br_0 wl_19 vdd gnd replica_cell_6t
Xrbc_20 bl_0 br_0 wl_20 vdd gnd replica_cell_6t
Xrbc_21 bl_0 br_0 wl_21 vdd gnd replica_cell_6t
Xrbc_22 bl_0 br_0 wl_22 vdd gnd replica_cell_6t
Xrbc_23 bl_0 br_0 wl_23 vdd gnd replica_cell_6t
Xrbc_24 bl_0 br_0 wl_24 vdd gnd replica_cell_6t
Xrbc_25 bl_0 br_0 wl_25 vdd gnd replica_cell_6t
Xrbc_26 bl_0 br_0 wl_26 vdd gnd replica_cell_6t
Xrbc_27 bl_0 br_0 wl_27 vdd gnd replica_cell_6t
Xrbc_28 bl_0 br_0 wl_28 vdd gnd replica_cell_6t
Xrbc_29 bl_0 br_0 wl_29 vdd gnd replica_cell_6t
Xrbc_30 bl_0 br_0 wl_30 vdd gnd replica_cell_6t
Xrbc_31 bl_0 br_0 wl_31 vdd gnd replica_cell_6t
Xrbc_32 bl_0 br_0 wl_32 vdd gnd replica_cell_6t
Xrbc_33 bl_0 br_0 wl_33 vdd gnd replica_cell_6t
Xrbc_34 bl_0 br_0 wl_34 vdd gnd replica_cell_6t
Xrbc_35 bl_0 br_0 wl_35 vdd gnd replica_cell_6t
Xrbc_36 bl_0 br_0 wl_36 vdd gnd replica_cell_6t
Xrbc_37 bl_0 br_0 wl_37 vdd gnd replica_cell_6t
Xrbc_38 bl_0 br_0 wl_38 vdd gnd replica_cell_6t
Xrbc_39 bl_0 br_0 wl_39 vdd gnd replica_cell_6t
Xrbc_40 bl_0 br_0 wl_40 vdd gnd replica_cell_6t
Xrbc_41 bl_0 br_0 wl_41 vdd gnd replica_cell_6t
Xrbc_42 bl_0 br_0 wl_42 vdd gnd replica_cell_6t
Xrbc_43 bl_0 br_0 wl_43 vdd gnd replica_cell_6t
Xrbc_44 bl_0 br_0 wl_44 vdd gnd replica_cell_6t
Xrbc_45 bl_0 br_0 wl_45 vdd gnd replica_cell_6t
Xrbc_46 bl_0 br_0 wl_46 vdd gnd replica_cell_6t
Xrbc_47 bl_0 br_0 wl_47 vdd gnd replica_cell_6t
Xrbc_48 bl_0 br_0 wl_48 vdd gnd replica_cell_6t
Xrbc_49 bl_0 br_0 wl_49 vdd gnd replica_cell_6t
Xrbc_50 bl_0 br_0 wl_50 vdd gnd replica_cell_6t
Xrbc_51 bl_0 br_0 wl_51 vdd gnd replica_cell_6t
Xrbc_52 bl_0 br_0 wl_52 vdd gnd replica_cell_6t
Xrbc_53 bl_0 br_0 wl_53 vdd gnd replica_cell_6t
Xrbc_54 bl_0 br_0 wl_54 vdd gnd replica_cell_6t
Xrbc_55 bl_0 br_0 wl_55 vdd gnd replica_cell_6t
Xrbc_56 bl_0 br_0 wl_56 vdd gnd replica_cell_6t
Xrbc_57 bl_0 br_0 wl_57 vdd gnd replica_cell_6t
Xrbc_58 bl_0 br_0 wl_58 vdd gnd replica_cell_6t
Xrbc_59 bl_0 br_0 wl_59 vdd gnd replica_cell_6t
Xrbc_60 bl_0 br_0 wl_60 vdd gnd replica_cell_6t
Xrbc_61 bl_0 br_0 wl_61 vdd gnd replica_cell_6t
Xrbc_62 bl_0 br_0 wl_62 vdd gnd replica_cell_6t
Xrbc_63 bl_0 br_0 wl_63 vdd gnd replica_cell_6t
Xrbc_64 bl_0 br_0 wl_64 vdd gnd replica_cell_6t
Xrbc_65 bl_0 br_0 wl_65 vdd gnd replica_cell_6t
Xrbc_66 bl_0 br_0 wl_66 vdd gnd replica_cell_6t
Xrbc_67 bl_0 br_0 wl_67 vdd gnd replica_cell_6t
Xrbc_68 bl_0 br_0 wl_68 vdd gnd replica_cell_6t
Xrbc_69 bl_0 br_0 wl_69 vdd gnd replica_cell_6t
Xrbc_70 bl_0 br_0 wl_70 vdd gnd replica_cell_6t
Xrbc_71 bl_0 br_0 wl_71 vdd gnd replica_cell_6t
Xrbc_72 bl_0 br_0 wl_72 vdd gnd replica_cell_6t
Xrbc_73 bl_0 br_0 wl_73 vdd gnd replica_cell_6t
Xrbc_74 bl_0 br_0 wl_74 vdd gnd replica_cell_6t
Xrbc_75 bl_0 br_0 wl_75 vdd gnd replica_cell_6t
Xrbc_76 bl_0 br_0 wl_76 vdd gnd replica_cell_6t
Xrbc_77 bl_0 br_0 wl_77 vdd gnd replica_cell_6t
Xrbc_78 bl_0 br_0 wl_78 vdd gnd replica_cell_6t
Xrbc_79 bl_0 br_0 wl_79 vdd gnd replica_cell_6t
Xrbc_80 bl_0 br_0 wl_80 vdd gnd replica_cell_6t
Xrbc_81 bl_0 br_0 wl_81 vdd gnd replica_cell_6t
Xrbc_82 bl_0 br_0 wl_82 vdd gnd replica_cell_6t
Xrbc_83 bl_0 br_0 wl_83 vdd gnd replica_cell_6t
Xrbc_84 bl_0 br_0 wl_84 vdd gnd replica_cell_6t
Xrbc_85 bl_0 br_0 wl_85 vdd gnd replica_cell_6t
Xrbc_86 bl_0 br_0 wl_86 vdd gnd replica_cell_6t
Xrbc_87 bl_0 br_0 wl_87 vdd gnd replica_cell_6t
Xrbc_88 bl_0 br_0 wl_88 vdd gnd replica_cell_6t
Xrbc_89 bl_0 br_0 wl_89 vdd gnd replica_cell_6t
Xrbc_90 bl_0 br_0 wl_90 vdd gnd replica_cell_6t
Xrbc_91 bl_0 br_0 wl_91 vdd gnd replica_cell_6t
Xrbc_92 bl_0 br_0 wl_92 vdd gnd replica_cell_6t
Xrbc_93 bl_0 br_0 wl_93 vdd gnd replica_cell_6t
Xrbc_94 bl_0 br_0 wl_94 vdd gnd replica_cell_6t
Xrbc_95 bl_0 br_0 wl_95 vdd gnd replica_cell_6t
Xrbc_96 bl_0 br_0 wl_96 vdd gnd replica_cell_6t
Xrbc_97 bl_0 br_0 wl_97 vdd gnd replica_cell_6t
Xrbc_98 bl_0 br_0 wl_98 vdd gnd replica_cell_6t
Xrbc_99 bl_0 br_0 wl_99 vdd gnd replica_cell_6t
Xrbc_100 bl_0 br_0 wl_100 vdd gnd replica_cell_6t
Xrbc_101 bl_0 br_0 wl_101 vdd gnd replica_cell_6t
Xrbc_102 bl_0 br_0 wl_102 vdd gnd replica_cell_6t
Xrbc_103 bl_0 br_0 wl_103 vdd gnd replica_cell_6t
Xrbc_104 bl_0 br_0 wl_104 vdd gnd replica_cell_6t
Xrbc_105 bl_0 br_0 wl_105 vdd gnd replica_cell_6t
Xrbc_106 bl_0 br_0 wl_106 vdd gnd replica_cell_6t
Xrbc_107 bl_0 br_0 wl_107 vdd gnd replica_cell_6t
Xrbc_108 bl_0 br_0 wl_108 vdd gnd replica_cell_6t
Xrbc_109 bl_0 br_0 wl_109 vdd gnd replica_cell_6t
Xrbc_110 bl_0 br_0 wl_110 vdd gnd replica_cell_6t
Xrbc_111 bl_0 br_0 wl_111 vdd gnd replica_cell_6t
Xrbc_112 bl_0 br_0 wl_112 vdd gnd replica_cell_6t
Xrbc_113 bl_0 br_0 wl_113 vdd gnd replica_cell_6t
Xrbc_114 bl_0 br_0 wl_114 vdd gnd replica_cell_6t
Xrbc_115 bl_0 br_0 wl_115 vdd gnd replica_cell_6t
Xrbc_116 bl_0 br_0 wl_116 vdd gnd replica_cell_6t
Xrbc_117 bl_0 br_0 wl_117 vdd gnd replica_cell_6t
Xrbc_118 bl_0 br_0 wl_118 vdd gnd replica_cell_6t
Xrbc_119 bl_0 br_0 wl_119 vdd gnd replica_cell_6t
Xrbc_120 bl_0 br_0 wl_120 vdd gnd replica_cell_6t
Xrbc_121 bl_0 br_0 wl_121 vdd gnd replica_cell_6t
Xrbc_122 bl_0 br_0 wl_122 vdd gnd replica_cell_6t
Xrbc_123 bl_0 br_0 wl_123 vdd gnd replica_cell_6t
Xrbc_124 bl_0 br_0 wl_124 vdd gnd replica_cell_6t
Xrbc_125 bl_0 br_0 wl_125 vdd gnd replica_cell_6t
Xrbc_126 bl_0 br_0 wl_126 vdd gnd replica_cell_6t
Xrbc_127 bl_0 br_0 wl_127 vdd gnd replica_cell_6t
Xrbc_128 bl_0 br_0 wl_128 vdd gnd replica_cell_6t
Xrbc_129 bl_0 br_0 wl_129 vdd gnd replica_cell_6t
Xrbc_130 bl_0 br_0 wl_130 vdd gnd dummy_cell_6t
.ENDS replica_column_0

.SUBCKT dummy_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* INPUT : wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 256
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c1 bl_1 br_1 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c2 bl_2 br_2 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c3 bl_3 br_3 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c4 bl_4 br_4 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c5 bl_5 br_5 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c6 bl_6 br_6 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c7 bl_7 br_7 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c8 bl_8 br_8 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c9 bl_9 br_9 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c10 bl_10 br_10 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c11 bl_11 br_11 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c12 bl_12 br_12 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c13 bl_13 br_13 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c14 bl_14 br_14 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c15 bl_15 br_15 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c16 bl_16 br_16 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c17 bl_17 br_17 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c18 bl_18 br_18 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c19 bl_19 br_19 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c20 bl_20 br_20 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c21 bl_21 br_21 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c22 bl_22 br_22 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c23 bl_23 br_23 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c24 bl_24 br_24 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c25 bl_25 br_25 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c26 bl_26 br_26 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c27 bl_27 br_27 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c28 bl_28 br_28 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c29 bl_29 br_29 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c30 bl_30 br_30 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c31 bl_31 br_31 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c32 bl_32 br_32 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c33 bl_33 br_33 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c34 bl_34 br_34 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c35 bl_35 br_35 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c36 bl_36 br_36 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c37 bl_37 br_37 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c38 bl_38 br_38 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c39 bl_39 br_39 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c40 bl_40 br_40 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c41 bl_41 br_41 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c42 bl_42 br_42 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c43 bl_43 br_43 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c44 bl_44 br_44 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c45 bl_45 br_45 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c46 bl_46 br_46 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c47 bl_47 br_47 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c48 bl_48 br_48 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c49 bl_49 br_49 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c50 bl_50 br_50 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c51 bl_51 br_51 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c52 bl_52 br_52 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c53 bl_53 br_53 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c54 bl_54 br_54 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c55 bl_55 br_55 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c56 bl_56 br_56 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c57 bl_57 br_57 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c58 bl_58 br_58 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c59 bl_59 br_59 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c60 bl_60 br_60 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c61 bl_61 br_61 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c62 bl_62 br_62 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c63 bl_63 br_63 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c64 bl_64 br_64 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c65 bl_65 br_65 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c66 bl_66 br_66 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c67 bl_67 br_67 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c68 bl_68 br_68 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c69 bl_69 br_69 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c70 bl_70 br_70 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c71 bl_71 br_71 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c72 bl_72 br_72 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c73 bl_73 br_73 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c74 bl_74 br_74 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c75 bl_75 br_75 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c76 bl_76 br_76 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c77 bl_77 br_77 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c78 bl_78 br_78 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c79 bl_79 br_79 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c80 bl_80 br_80 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c81 bl_81 br_81 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c82 bl_82 br_82 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c83 bl_83 br_83 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c84 bl_84 br_84 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c85 bl_85 br_85 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c86 bl_86 br_86 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c87 bl_87 br_87 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c88 bl_88 br_88 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c89 bl_89 br_89 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c90 bl_90 br_90 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c91 bl_91 br_91 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c92 bl_92 br_92 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c93 bl_93 br_93 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c94 bl_94 br_94 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c95 bl_95 br_95 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c96 bl_96 br_96 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c97 bl_97 br_97 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c98 bl_98 br_98 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c99 bl_99 br_99 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c100 bl_100 br_100 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c101 bl_101 br_101 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c102 bl_102 br_102 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c103 bl_103 br_103 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c104 bl_104 br_104 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c105 bl_105 br_105 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c106 bl_106 br_106 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c107 bl_107 br_107 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c108 bl_108 br_108 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c109 bl_109 br_109 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c110 bl_110 br_110 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c111 bl_111 br_111 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c112 bl_112 br_112 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c113 bl_113 br_113 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c114 bl_114 br_114 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c115 bl_115 br_115 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c116 bl_116 br_116 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c117 bl_117 br_117 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c118 bl_118 br_118 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c119 bl_119 br_119 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c120 bl_120 br_120 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c121 bl_121 br_121 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c122 bl_122 br_122 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c123 bl_123 br_123 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c124 bl_124 br_124 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c125 bl_125 br_125 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c126 bl_126 br_126 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c127 bl_127 br_127 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c128 bl_128 br_128 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c129 bl_129 br_129 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c130 bl_130 br_130 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c131 bl_131 br_131 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c132 bl_132 br_132 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c133 bl_133 br_133 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c134 bl_134 br_134 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c135 bl_135 br_135 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c136 bl_136 br_136 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c137 bl_137 br_137 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c138 bl_138 br_138 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c139 bl_139 br_139 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c140 bl_140 br_140 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c141 bl_141 br_141 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c142 bl_142 br_142 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c143 bl_143 br_143 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c144 bl_144 br_144 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c145 bl_145 br_145 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c146 bl_146 br_146 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c147 bl_147 br_147 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c148 bl_148 br_148 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c149 bl_149 br_149 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c150 bl_150 br_150 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c151 bl_151 br_151 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c152 bl_152 br_152 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c153 bl_153 br_153 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c154 bl_154 br_154 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c155 bl_155 br_155 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c156 bl_156 br_156 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c157 bl_157 br_157 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c158 bl_158 br_158 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c159 bl_159 br_159 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c160 bl_160 br_160 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c161 bl_161 br_161 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c162 bl_162 br_162 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c163 bl_163 br_163 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c164 bl_164 br_164 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c165 bl_165 br_165 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c166 bl_166 br_166 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c167 bl_167 br_167 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c168 bl_168 br_168 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c169 bl_169 br_169 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c170 bl_170 br_170 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c171 bl_171 br_171 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c172 bl_172 br_172 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c173 bl_173 br_173 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c174 bl_174 br_174 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c175 bl_175 br_175 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c176 bl_176 br_176 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c177 bl_177 br_177 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c178 bl_178 br_178 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c179 bl_179 br_179 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c180 bl_180 br_180 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c181 bl_181 br_181 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c182 bl_182 br_182 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c183 bl_183 br_183 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c184 bl_184 br_184 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c185 bl_185 br_185 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c186 bl_186 br_186 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c187 bl_187 br_187 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c188 bl_188 br_188 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c189 bl_189 br_189 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c190 bl_190 br_190 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c191 bl_191 br_191 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c192 bl_192 br_192 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c193 bl_193 br_193 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c194 bl_194 br_194 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c195 bl_195 br_195 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c196 bl_196 br_196 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c197 bl_197 br_197 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c198 bl_198 br_198 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c199 bl_199 br_199 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c200 bl_200 br_200 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c201 bl_201 br_201 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c202 bl_202 br_202 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c203 bl_203 br_203 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c204 bl_204 br_204 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c205 bl_205 br_205 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c206 bl_206 br_206 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c207 bl_207 br_207 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c208 bl_208 br_208 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c209 bl_209 br_209 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c210 bl_210 br_210 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c211 bl_211 br_211 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c212 bl_212 br_212 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c213 bl_213 br_213 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c214 bl_214 br_214 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c215 bl_215 br_215 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c216 bl_216 br_216 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c217 bl_217 br_217 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c218 bl_218 br_218 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c219 bl_219 br_219 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c220 bl_220 br_220 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c221 bl_221 br_221 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c222 bl_222 br_222 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c223 bl_223 br_223 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c224 bl_224 br_224 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c225 bl_225 br_225 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c226 bl_226 br_226 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c227 bl_227 br_227 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c228 bl_228 br_228 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c229 bl_229 br_229 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c230 bl_230 br_230 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c231 bl_231 br_231 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c232 bl_232 br_232 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c233 bl_233 br_233 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c234 bl_234 br_234 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c235 bl_235 br_235 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c236 bl_236 br_236 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c237 bl_237 br_237 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c238 bl_238 br_238 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c239 bl_239 br_239 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c240 bl_240 br_240 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c241 bl_241 br_241 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c242 bl_242 br_242 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c243 bl_243 br_243 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c244 bl_244 br_244 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c245 bl_245 br_245 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c246 bl_246 br_246 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c247 bl_247 br_247 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c248 bl_248 br_248 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c249 bl_249 br_249 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c250 bl_250 br_250 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c251 bl_251 br_251 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c252 bl_252 br_252 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c253 bl_253 br_253 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c254 bl_254 br_254 wl_0 vdd gnd dummy_cell_6t
Xbit_r0_c255 bl_255 br_255 wl_0 vdd gnd dummy_cell_6t
.ENDS dummy_array_0

.SUBCKT dummy_array_1 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* POWER : vdd 
* GROUND: gnd 
* rows: 131 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd dummy_cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd dummy_cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd dummy_cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd dummy_cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd dummy_cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd dummy_cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd dummy_cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd dummy_cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd dummy_cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd dummy_cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd dummy_cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd dummy_cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd dummy_cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd dummy_cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd dummy_cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd dummy_cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd dummy_cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd dummy_cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd dummy_cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd dummy_cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd dummy_cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd dummy_cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd dummy_cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd dummy_cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd dummy_cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd dummy_cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd dummy_cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd dummy_cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd dummy_cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd dummy_cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd dummy_cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd dummy_cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd dummy_cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd dummy_cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd dummy_cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd dummy_cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd dummy_cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd dummy_cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd dummy_cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd dummy_cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd dummy_cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd dummy_cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd dummy_cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd dummy_cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd dummy_cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd dummy_cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd dummy_cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd dummy_cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd dummy_cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd dummy_cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd dummy_cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd dummy_cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd dummy_cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd dummy_cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd dummy_cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd dummy_cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd dummy_cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd dummy_cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd dummy_cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd dummy_cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd dummy_cell_6t
Xbit_r128_c0 bl_0 br_0 wl_128 vdd gnd dummy_cell_6t
Xbit_r129_c0 bl_0 br_0 wl_129 vdd gnd dummy_cell_6t
Xbit_r130_c0 bl_0 br_0 wl_130 vdd gnd dummy_cell_6t
.ENDS dummy_array_1

.SUBCKT dummy_array_2 bl_0 br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_128 wl_129 wl_130 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : wl_128 
* INPUT : wl_129 
* INPUT : wl_130 
* POWER : vdd 
* GROUND: gnd 
* rows: 131 cols: 1
Xbit_r0_c0 bl_0 br_0 wl_0 vdd gnd dummy_cell_6t
Xbit_r1_c0 bl_0 br_0 wl_1 vdd gnd dummy_cell_6t
Xbit_r2_c0 bl_0 br_0 wl_2 vdd gnd dummy_cell_6t
Xbit_r3_c0 bl_0 br_0 wl_3 vdd gnd dummy_cell_6t
Xbit_r4_c0 bl_0 br_0 wl_4 vdd gnd dummy_cell_6t
Xbit_r5_c0 bl_0 br_0 wl_5 vdd gnd dummy_cell_6t
Xbit_r6_c0 bl_0 br_0 wl_6 vdd gnd dummy_cell_6t
Xbit_r7_c0 bl_0 br_0 wl_7 vdd gnd dummy_cell_6t
Xbit_r8_c0 bl_0 br_0 wl_8 vdd gnd dummy_cell_6t
Xbit_r9_c0 bl_0 br_0 wl_9 vdd gnd dummy_cell_6t
Xbit_r10_c0 bl_0 br_0 wl_10 vdd gnd dummy_cell_6t
Xbit_r11_c0 bl_0 br_0 wl_11 vdd gnd dummy_cell_6t
Xbit_r12_c0 bl_0 br_0 wl_12 vdd gnd dummy_cell_6t
Xbit_r13_c0 bl_0 br_0 wl_13 vdd gnd dummy_cell_6t
Xbit_r14_c0 bl_0 br_0 wl_14 vdd gnd dummy_cell_6t
Xbit_r15_c0 bl_0 br_0 wl_15 vdd gnd dummy_cell_6t
Xbit_r16_c0 bl_0 br_0 wl_16 vdd gnd dummy_cell_6t
Xbit_r17_c0 bl_0 br_0 wl_17 vdd gnd dummy_cell_6t
Xbit_r18_c0 bl_0 br_0 wl_18 vdd gnd dummy_cell_6t
Xbit_r19_c0 bl_0 br_0 wl_19 vdd gnd dummy_cell_6t
Xbit_r20_c0 bl_0 br_0 wl_20 vdd gnd dummy_cell_6t
Xbit_r21_c0 bl_0 br_0 wl_21 vdd gnd dummy_cell_6t
Xbit_r22_c0 bl_0 br_0 wl_22 vdd gnd dummy_cell_6t
Xbit_r23_c0 bl_0 br_0 wl_23 vdd gnd dummy_cell_6t
Xbit_r24_c0 bl_0 br_0 wl_24 vdd gnd dummy_cell_6t
Xbit_r25_c0 bl_0 br_0 wl_25 vdd gnd dummy_cell_6t
Xbit_r26_c0 bl_0 br_0 wl_26 vdd gnd dummy_cell_6t
Xbit_r27_c0 bl_0 br_0 wl_27 vdd gnd dummy_cell_6t
Xbit_r28_c0 bl_0 br_0 wl_28 vdd gnd dummy_cell_6t
Xbit_r29_c0 bl_0 br_0 wl_29 vdd gnd dummy_cell_6t
Xbit_r30_c0 bl_0 br_0 wl_30 vdd gnd dummy_cell_6t
Xbit_r31_c0 bl_0 br_0 wl_31 vdd gnd dummy_cell_6t
Xbit_r32_c0 bl_0 br_0 wl_32 vdd gnd dummy_cell_6t
Xbit_r33_c0 bl_0 br_0 wl_33 vdd gnd dummy_cell_6t
Xbit_r34_c0 bl_0 br_0 wl_34 vdd gnd dummy_cell_6t
Xbit_r35_c0 bl_0 br_0 wl_35 vdd gnd dummy_cell_6t
Xbit_r36_c0 bl_0 br_0 wl_36 vdd gnd dummy_cell_6t
Xbit_r37_c0 bl_0 br_0 wl_37 vdd gnd dummy_cell_6t
Xbit_r38_c0 bl_0 br_0 wl_38 vdd gnd dummy_cell_6t
Xbit_r39_c0 bl_0 br_0 wl_39 vdd gnd dummy_cell_6t
Xbit_r40_c0 bl_0 br_0 wl_40 vdd gnd dummy_cell_6t
Xbit_r41_c0 bl_0 br_0 wl_41 vdd gnd dummy_cell_6t
Xbit_r42_c0 bl_0 br_0 wl_42 vdd gnd dummy_cell_6t
Xbit_r43_c0 bl_0 br_0 wl_43 vdd gnd dummy_cell_6t
Xbit_r44_c0 bl_0 br_0 wl_44 vdd gnd dummy_cell_6t
Xbit_r45_c0 bl_0 br_0 wl_45 vdd gnd dummy_cell_6t
Xbit_r46_c0 bl_0 br_0 wl_46 vdd gnd dummy_cell_6t
Xbit_r47_c0 bl_0 br_0 wl_47 vdd gnd dummy_cell_6t
Xbit_r48_c0 bl_0 br_0 wl_48 vdd gnd dummy_cell_6t
Xbit_r49_c0 bl_0 br_0 wl_49 vdd gnd dummy_cell_6t
Xbit_r50_c0 bl_0 br_0 wl_50 vdd gnd dummy_cell_6t
Xbit_r51_c0 bl_0 br_0 wl_51 vdd gnd dummy_cell_6t
Xbit_r52_c0 bl_0 br_0 wl_52 vdd gnd dummy_cell_6t
Xbit_r53_c0 bl_0 br_0 wl_53 vdd gnd dummy_cell_6t
Xbit_r54_c0 bl_0 br_0 wl_54 vdd gnd dummy_cell_6t
Xbit_r55_c0 bl_0 br_0 wl_55 vdd gnd dummy_cell_6t
Xbit_r56_c0 bl_0 br_0 wl_56 vdd gnd dummy_cell_6t
Xbit_r57_c0 bl_0 br_0 wl_57 vdd gnd dummy_cell_6t
Xbit_r58_c0 bl_0 br_0 wl_58 vdd gnd dummy_cell_6t
Xbit_r59_c0 bl_0 br_0 wl_59 vdd gnd dummy_cell_6t
Xbit_r60_c0 bl_0 br_0 wl_60 vdd gnd dummy_cell_6t
Xbit_r61_c0 bl_0 br_0 wl_61 vdd gnd dummy_cell_6t
Xbit_r62_c0 bl_0 br_0 wl_62 vdd gnd dummy_cell_6t
Xbit_r63_c0 bl_0 br_0 wl_63 vdd gnd dummy_cell_6t
Xbit_r64_c0 bl_0 br_0 wl_64 vdd gnd dummy_cell_6t
Xbit_r65_c0 bl_0 br_0 wl_65 vdd gnd dummy_cell_6t
Xbit_r66_c0 bl_0 br_0 wl_66 vdd gnd dummy_cell_6t
Xbit_r67_c0 bl_0 br_0 wl_67 vdd gnd dummy_cell_6t
Xbit_r68_c0 bl_0 br_0 wl_68 vdd gnd dummy_cell_6t
Xbit_r69_c0 bl_0 br_0 wl_69 vdd gnd dummy_cell_6t
Xbit_r70_c0 bl_0 br_0 wl_70 vdd gnd dummy_cell_6t
Xbit_r71_c0 bl_0 br_0 wl_71 vdd gnd dummy_cell_6t
Xbit_r72_c0 bl_0 br_0 wl_72 vdd gnd dummy_cell_6t
Xbit_r73_c0 bl_0 br_0 wl_73 vdd gnd dummy_cell_6t
Xbit_r74_c0 bl_0 br_0 wl_74 vdd gnd dummy_cell_6t
Xbit_r75_c0 bl_0 br_0 wl_75 vdd gnd dummy_cell_6t
Xbit_r76_c0 bl_0 br_0 wl_76 vdd gnd dummy_cell_6t
Xbit_r77_c0 bl_0 br_0 wl_77 vdd gnd dummy_cell_6t
Xbit_r78_c0 bl_0 br_0 wl_78 vdd gnd dummy_cell_6t
Xbit_r79_c0 bl_0 br_0 wl_79 vdd gnd dummy_cell_6t
Xbit_r80_c0 bl_0 br_0 wl_80 vdd gnd dummy_cell_6t
Xbit_r81_c0 bl_0 br_0 wl_81 vdd gnd dummy_cell_6t
Xbit_r82_c0 bl_0 br_0 wl_82 vdd gnd dummy_cell_6t
Xbit_r83_c0 bl_0 br_0 wl_83 vdd gnd dummy_cell_6t
Xbit_r84_c0 bl_0 br_0 wl_84 vdd gnd dummy_cell_6t
Xbit_r85_c0 bl_0 br_0 wl_85 vdd gnd dummy_cell_6t
Xbit_r86_c0 bl_0 br_0 wl_86 vdd gnd dummy_cell_6t
Xbit_r87_c0 bl_0 br_0 wl_87 vdd gnd dummy_cell_6t
Xbit_r88_c0 bl_0 br_0 wl_88 vdd gnd dummy_cell_6t
Xbit_r89_c0 bl_0 br_0 wl_89 vdd gnd dummy_cell_6t
Xbit_r90_c0 bl_0 br_0 wl_90 vdd gnd dummy_cell_6t
Xbit_r91_c0 bl_0 br_0 wl_91 vdd gnd dummy_cell_6t
Xbit_r92_c0 bl_0 br_0 wl_92 vdd gnd dummy_cell_6t
Xbit_r93_c0 bl_0 br_0 wl_93 vdd gnd dummy_cell_6t
Xbit_r94_c0 bl_0 br_0 wl_94 vdd gnd dummy_cell_6t
Xbit_r95_c0 bl_0 br_0 wl_95 vdd gnd dummy_cell_6t
Xbit_r96_c0 bl_0 br_0 wl_96 vdd gnd dummy_cell_6t
Xbit_r97_c0 bl_0 br_0 wl_97 vdd gnd dummy_cell_6t
Xbit_r98_c0 bl_0 br_0 wl_98 vdd gnd dummy_cell_6t
Xbit_r99_c0 bl_0 br_0 wl_99 vdd gnd dummy_cell_6t
Xbit_r100_c0 bl_0 br_0 wl_100 vdd gnd dummy_cell_6t
Xbit_r101_c0 bl_0 br_0 wl_101 vdd gnd dummy_cell_6t
Xbit_r102_c0 bl_0 br_0 wl_102 vdd gnd dummy_cell_6t
Xbit_r103_c0 bl_0 br_0 wl_103 vdd gnd dummy_cell_6t
Xbit_r104_c0 bl_0 br_0 wl_104 vdd gnd dummy_cell_6t
Xbit_r105_c0 bl_0 br_0 wl_105 vdd gnd dummy_cell_6t
Xbit_r106_c0 bl_0 br_0 wl_106 vdd gnd dummy_cell_6t
Xbit_r107_c0 bl_0 br_0 wl_107 vdd gnd dummy_cell_6t
Xbit_r108_c0 bl_0 br_0 wl_108 vdd gnd dummy_cell_6t
Xbit_r109_c0 bl_0 br_0 wl_109 vdd gnd dummy_cell_6t
Xbit_r110_c0 bl_0 br_0 wl_110 vdd gnd dummy_cell_6t
Xbit_r111_c0 bl_0 br_0 wl_111 vdd gnd dummy_cell_6t
Xbit_r112_c0 bl_0 br_0 wl_112 vdd gnd dummy_cell_6t
Xbit_r113_c0 bl_0 br_0 wl_113 vdd gnd dummy_cell_6t
Xbit_r114_c0 bl_0 br_0 wl_114 vdd gnd dummy_cell_6t
Xbit_r115_c0 bl_0 br_0 wl_115 vdd gnd dummy_cell_6t
Xbit_r116_c0 bl_0 br_0 wl_116 vdd gnd dummy_cell_6t
Xbit_r117_c0 bl_0 br_0 wl_117 vdd gnd dummy_cell_6t
Xbit_r118_c0 bl_0 br_0 wl_118 vdd gnd dummy_cell_6t
Xbit_r119_c0 bl_0 br_0 wl_119 vdd gnd dummy_cell_6t
Xbit_r120_c0 bl_0 br_0 wl_120 vdd gnd dummy_cell_6t
Xbit_r121_c0 bl_0 br_0 wl_121 vdd gnd dummy_cell_6t
Xbit_r122_c0 bl_0 br_0 wl_122 vdd gnd dummy_cell_6t
Xbit_r123_c0 bl_0 br_0 wl_123 vdd gnd dummy_cell_6t
Xbit_r124_c0 bl_0 br_0 wl_124 vdd gnd dummy_cell_6t
Xbit_r125_c0 bl_0 br_0 wl_125 vdd gnd dummy_cell_6t
Xbit_r126_c0 bl_0 br_0 wl_126 vdd gnd dummy_cell_6t
Xbit_r127_c0 bl_0 br_0 wl_127 vdd gnd dummy_cell_6t
Xbit_r128_c0 bl_0 br_0 wl_128 vdd gnd dummy_cell_6t
Xbit_r129_c0 bl_0 br_0 wl_129 vdd gnd dummy_cell_6t
Xbit_r130_c0 bl_0 br_0 wl_130 vdd gnd dummy_cell_6t
.ENDS dummy_array_2

.SUBCKT replica_bitcell_array_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 rbl_wl_0 vdd gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : bl_64 
* INOUT : br_64 
* INOUT : bl_65 
* INOUT : br_65 
* INOUT : bl_66 
* INOUT : br_66 
* INOUT : bl_67 
* INOUT : br_67 
* INOUT : bl_68 
* INOUT : br_68 
* INOUT : bl_69 
* INOUT : br_69 
* INOUT : bl_70 
* INOUT : br_70 
* INOUT : bl_71 
* INOUT : br_71 
* INOUT : bl_72 
* INOUT : br_72 
* INOUT : bl_73 
* INOUT : br_73 
* INOUT : bl_74 
* INOUT : br_74 
* INOUT : bl_75 
* INOUT : br_75 
* INOUT : bl_76 
* INOUT : br_76 
* INOUT : bl_77 
* INOUT : br_77 
* INOUT : bl_78 
* INOUT : br_78 
* INOUT : bl_79 
* INOUT : br_79 
* INOUT : bl_80 
* INOUT : br_80 
* INOUT : bl_81 
* INOUT : br_81 
* INOUT : bl_82 
* INOUT : br_82 
* INOUT : bl_83 
* INOUT : br_83 
* INOUT : bl_84 
* INOUT : br_84 
* INOUT : bl_85 
* INOUT : br_85 
* INOUT : bl_86 
* INOUT : br_86 
* INOUT : bl_87 
* INOUT : br_87 
* INOUT : bl_88 
* INOUT : br_88 
* INOUT : bl_89 
* INOUT : br_89 
* INOUT : bl_90 
* INOUT : br_90 
* INOUT : bl_91 
* INOUT : br_91 
* INOUT : bl_92 
* INOUT : br_92 
* INOUT : bl_93 
* INOUT : br_93 
* INOUT : bl_94 
* INOUT : br_94 
* INOUT : bl_95 
* INOUT : br_95 
* INOUT : bl_96 
* INOUT : br_96 
* INOUT : bl_97 
* INOUT : br_97 
* INOUT : bl_98 
* INOUT : br_98 
* INOUT : bl_99 
* INOUT : br_99 
* INOUT : bl_100 
* INOUT : br_100 
* INOUT : bl_101 
* INOUT : br_101 
* INOUT : bl_102 
* INOUT : br_102 
* INOUT : bl_103 
* INOUT : br_103 
* INOUT : bl_104 
* INOUT : br_104 
* INOUT : bl_105 
* INOUT : br_105 
* INOUT : bl_106 
* INOUT : br_106 
* INOUT : bl_107 
* INOUT : br_107 
* INOUT : bl_108 
* INOUT : br_108 
* INOUT : bl_109 
* INOUT : br_109 
* INOUT : bl_110 
* INOUT : br_110 
* INOUT : bl_111 
* INOUT : br_111 
* INOUT : bl_112 
* INOUT : br_112 
* INOUT : bl_113 
* INOUT : br_113 
* INOUT : bl_114 
* INOUT : br_114 
* INOUT : bl_115 
* INOUT : br_115 
* INOUT : bl_116 
* INOUT : br_116 
* INOUT : bl_117 
* INOUT : br_117 
* INOUT : bl_118 
* INOUT : br_118 
* INOUT : bl_119 
* INOUT : br_119 
* INOUT : bl_120 
* INOUT : br_120 
* INOUT : bl_121 
* INOUT : br_121 
* INOUT : bl_122 
* INOUT : br_122 
* INOUT : bl_123 
* INOUT : br_123 
* INOUT : bl_124 
* INOUT : br_124 
* INOUT : bl_125 
* INOUT : br_125 
* INOUT : bl_126 
* INOUT : br_126 
* INOUT : bl_127 
* INOUT : br_127 
* INOUT : bl_128 
* INOUT : br_128 
* INOUT : bl_129 
* INOUT : br_129 
* INOUT : bl_130 
* INOUT : br_130 
* INOUT : bl_131 
* INOUT : br_131 
* INOUT : bl_132 
* INOUT : br_132 
* INOUT : bl_133 
* INOUT : br_133 
* INOUT : bl_134 
* INOUT : br_134 
* INOUT : bl_135 
* INOUT : br_135 
* INOUT : bl_136 
* INOUT : br_136 
* INOUT : bl_137 
* INOUT : br_137 
* INOUT : bl_138 
* INOUT : br_138 
* INOUT : bl_139 
* INOUT : br_139 
* INOUT : bl_140 
* INOUT : br_140 
* INOUT : bl_141 
* INOUT : br_141 
* INOUT : bl_142 
* INOUT : br_142 
* INOUT : bl_143 
* INOUT : br_143 
* INOUT : bl_144 
* INOUT : br_144 
* INOUT : bl_145 
* INOUT : br_145 
* INOUT : bl_146 
* INOUT : br_146 
* INOUT : bl_147 
* INOUT : br_147 
* INOUT : bl_148 
* INOUT : br_148 
* INOUT : bl_149 
* INOUT : br_149 
* INOUT : bl_150 
* INOUT : br_150 
* INOUT : bl_151 
* INOUT : br_151 
* INOUT : bl_152 
* INOUT : br_152 
* INOUT : bl_153 
* INOUT : br_153 
* INOUT : bl_154 
* INOUT : br_154 
* INOUT : bl_155 
* INOUT : br_155 
* INOUT : bl_156 
* INOUT : br_156 
* INOUT : bl_157 
* INOUT : br_157 
* INOUT : bl_158 
* INOUT : br_158 
* INOUT : bl_159 
* INOUT : br_159 
* INOUT : bl_160 
* INOUT : br_160 
* INOUT : bl_161 
* INOUT : br_161 
* INOUT : bl_162 
* INOUT : br_162 
* INOUT : bl_163 
* INOUT : br_163 
* INOUT : bl_164 
* INOUT : br_164 
* INOUT : bl_165 
* INOUT : br_165 
* INOUT : bl_166 
* INOUT : br_166 
* INOUT : bl_167 
* INOUT : br_167 
* INOUT : bl_168 
* INOUT : br_168 
* INOUT : bl_169 
* INOUT : br_169 
* INOUT : bl_170 
* INOUT : br_170 
* INOUT : bl_171 
* INOUT : br_171 
* INOUT : bl_172 
* INOUT : br_172 
* INOUT : bl_173 
* INOUT : br_173 
* INOUT : bl_174 
* INOUT : br_174 
* INOUT : bl_175 
* INOUT : br_175 
* INOUT : bl_176 
* INOUT : br_176 
* INOUT : bl_177 
* INOUT : br_177 
* INOUT : bl_178 
* INOUT : br_178 
* INOUT : bl_179 
* INOUT : br_179 
* INOUT : bl_180 
* INOUT : br_180 
* INOUT : bl_181 
* INOUT : br_181 
* INOUT : bl_182 
* INOUT : br_182 
* INOUT : bl_183 
* INOUT : br_183 
* INOUT : bl_184 
* INOUT : br_184 
* INOUT : bl_185 
* INOUT : br_185 
* INOUT : bl_186 
* INOUT : br_186 
* INOUT : bl_187 
* INOUT : br_187 
* INOUT : bl_188 
* INOUT : br_188 
* INOUT : bl_189 
* INOUT : br_189 
* INOUT : bl_190 
* INOUT : br_190 
* INOUT : bl_191 
* INOUT : br_191 
* INOUT : bl_192 
* INOUT : br_192 
* INOUT : bl_193 
* INOUT : br_193 
* INOUT : bl_194 
* INOUT : br_194 
* INOUT : bl_195 
* INOUT : br_195 
* INOUT : bl_196 
* INOUT : br_196 
* INOUT : bl_197 
* INOUT : br_197 
* INOUT : bl_198 
* INOUT : br_198 
* INOUT : bl_199 
* INOUT : br_199 
* INOUT : bl_200 
* INOUT : br_200 
* INOUT : bl_201 
* INOUT : br_201 
* INOUT : bl_202 
* INOUT : br_202 
* INOUT : bl_203 
* INOUT : br_203 
* INOUT : bl_204 
* INOUT : br_204 
* INOUT : bl_205 
* INOUT : br_205 
* INOUT : bl_206 
* INOUT : br_206 
* INOUT : bl_207 
* INOUT : br_207 
* INOUT : bl_208 
* INOUT : br_208 
* INOUT : bl_209 
* INOUT : br_209 
* INOUT : bl_210 
* INOUT : br_210 
* INOUT : bl_211 
* INOUT : br_211 
* INOUT : bl_212 
* INOUT : br_212 
* INOUT : bl_213 
* INOUT : br_213 
* INOUT : bl_214 
* INOUT : br_214 
* INOUT : bl_215 
* INOUT : br_215 
* INOUT : bl_216 
* INOUT : br_216 
* INOUT : bl_217 
* INOUT : br_217 
* INOUT : bl_218 
* INOUT : br_218 
* INOUT : bl_219 
* INOUT : br_219 
* INOUT : bl_220 
* INOUT : br_220 
* INOUT : bl_221 
* INOUT : br_221 
* INOUT : bl_222 
* INOUT : br_222 
* INOUT : bl_223 
* INOUT : br_223 
* INOUT : bl_224 
* INOUT : br_224 
* INOUT : bl_225 
* INOUT : br_225 
* INOUT : bl_226 
* INOUT : br_226 
* INOUT : bl_227 
* INOUT : br_227 
* INOUT : bl_228 
* INOUT : br_228 
* INOUT : bl_229 
* INOUT : br_229 
* INOUT : bl_230 
* INOUT : br_230 
* INOUT : bl_231 
* INOUT : br_231 
* INOUT : bl_232 
* INOUT : br_232 
* INOUT : bl_233 
* INOUT : br_233 
* INOUT : bl_234 
* INOUT : br_234 
* INOUT : bl_235 
* INOUT : br_235 
* INOUT : bl_236 
* INOUT : br_236 
* INOUT : bl_237 
* INOUT : br_237 
* INOUT : bl_238 
* INOUT : br_238 
* INOUT : bl_239 
* INOUT : br_239 
* INOUT : bl_240 
* INOUT : br_240 
* INOUT : bl_241 
* INOUT : br_241 
* INOUT : bl_242 
* INOUT : br_242 
* INOUT : bl_243 
* INOUT : br_243 
* INOUT : bl_244 
* INOUT : br_244 
* INOUT : bl_245 
* INOUT : br_245 
* INOUT : bl_246 
* INOUT : br_246 
* INOUT : bl_247 
* INOUT : br_247 
* INOUT : bl_248 
* INOUT : br_248 
* INOUT : bl_249 
* INOUT : br_249 
* INOUT : bl_250 
* INOUT : br_250 
* INOUT : bl_251 
* INOUT : br_251 
* INOUT : bl_252 
* INOUT : br_252 
* INOUT : bl_253 
* INOUT : br_253 
* INOUT : bl_254 
* INOUT : br_254 
* INOUT : bl_255 
* INOUT : br_255 
* OUTPUT: rbl_bl_0 
* OUTPUT: rbl_br_0 
* INPUT : wl_0 
* INPUT : wl_1 
* INPUT : wl_2 
* INPUT : wl_3 
* INPUT : wl_4 
* INPUT : wl_5 
* INPUT : wl_6 
* INPUT : wl_7 
* INPUT : wl_8 
* INPUT : wl_9 
* INPUT : wl_10 
* INPUT : wl_11 
* INPUT : wl_12 
* INPUT : wl_13 
* INPUT : wl_14 
* INPUT : wl_15 
* INPUT : wl_16 
* INPUT : wl_17 
* INPUT : wl_18 
* INPUT : wl_19 
* INPUT : wl_20 
* INPUT : wl_21 
* INPUT : wl_22 
* INPUT : wl_23 
* INPUT : wl_24 
* INPUT : wl_25 
* INPUT : wl_26 
* INPUT : wl_27 
* INPUT : wl_28 
* INPUT : wl_29 
* INPUT : wl_30 
* INPUT : wl_31 
* INPUT : wl_32 
* INPUT : wl_33 
* INPUT : wl_34 
* INPUT : wl_35 
* INPUT : wl_36 
* INPUT : wl_37 
* INPUT : wl_38 
* INPUT : wl_39 
* INPUT : wl_40 
* INPUT : wl_41 
* INPUT : wl_42 
* INPUT : wl_43 
* INPUT : wl_44 
* INPUT : wl_45 
* INPUT : wl_46 
* INPUT : wl_47 
* INPUT : wl_48 
* INPUT : wl_49 
* INPUT : wl_50 
* INPUT : wl_51 
* INPUT : wl_52 
* INPUT : wl_53 
* INPUT : wl_54 
* INPUT : wl_55 
* INPUT : wl_56 
* INPUT : wl_57 
* INPUT : wl_58 
* INPUT : wl_59 
* INPUT : wl_60 
* INPUT : wl_61 
* INPUT : wl_62 
* INPUT : wl_63 
* INPUT : wl_64 
* INPUT : wl_65 
* INPUT : wl_66 
* INPUT : wl_67 
* INPUT : wl_68 
* INPUT : wl_69 
* INPUT : wl_70 
* INPUT : wl_71 
* INPUT : wl_72 
* INPUT : wl_73 
* INPUT : wl_74 
* INPUT : wl_75 
* INPUT : wl_76 
* INPUT : wl_77 
* INPUT : wl_78 
* INPUT : wl_79 
* INPUT : wl_80 
* INPUT : wl_81 
* INPUT : wl_82 
* INPUT : wl_83 
* INPUT : wl_84 
* INPUT : wl_85 
* INPUT : wl_86 
* INPUT : wl_87 
* INPUT : wl_88 
* INPUT : wl_89 
* INPUT : wl_90 
* INPUT : wl_91 
* INPUT : wl_92 
* INPUT : wl_93 
* INPUT : wl_94 
* INPUT : wl_95 
* INPUT : wl_96 
* INPUT : wl_97 
* INPUT : wl_98 
* INPUT : wl_99 
* INPUT : wl_100 
* INPUT : wl_101 
* INPUT : wl_102 
* INPUT : wl_103 
* INPUT : wl_104 
* INPUT : wl_105 
* INPUT : wl_106 
* INPUT : wl_107 
* INPUT : wl_108 
* INPUT : wl_109 
* INPUT : wl_110 
* INPUT : wl_111 
* INPUT : wl_112 
* INPUT : wl_113 
* INPUT : wl_114 
* INPUT : wl_115 
* INPUT : wl_116 
* INPUT : wl_117 
* INPUT : wl_118 
* INPUT : wl_119 
* INPUT : wl_120 
* INPUT : wl_121 
* INPUT : wl_122 
* INPUT : wl_123 
* INPUT : wl_124 
* INPUT : wl_125 
* INPUT : wl_126 
* INPUT : wl_127 
* INPUT : rbl_wl_0 
* POWER : vdd 
* GROUND: gnd 
* rows: 128 cols: 256
Xbitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 vdd gnd bitcell_array_0
Xreplica_col_0 rbl_bl_0 rbl_br_0 dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 dummy_wl_top vdd gnd replica_column_0
Xdummy_row_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_wl_0 vdd gnd dummy_array_0
Xdummy_row_bot bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_bot vdd gnd dummy_array_0
Xdummy_row_top bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dummy_wl_top vdd gnd dummy_array_0
Xdummy_col_left dummy_bl_left dummy_br_left dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 dummy_wl_top vdd gnd dummy_array_1
Xdummy_col_right dummy_bl_right dummy_br_right dummy_wl_bot rbl_wl_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 dummy_wl_top vdd gnd dummy_array_2
.ENDS replica_bitcell_array_0

.SUBCKT pinv_6 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_6

.SUBCKT pnand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand3_1

.SUBCKT hierarchical_predecode3x8_1 in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0 in_0 inbar_0 vdd gnd pinv_6
Xpre_inv_1 in_1 inbar_1 vdd gnd pinv_6
Xpre_inv_2 in_2 inbar_2 vdd gnd pinv_6
Xpre_nand_inv_0 Z_0 out_0 vdd gnd pinv_6
Xpre_nand_inv_1 Z_1 out_1 vdd gnd pinv_6
Xpre_nand_inv_2 Z_2 out_2 vdd gnd pinv_6
Xpre_nand_inv_3 Z_3 out_3 vdd gnd pinv_6
Xpre_nand_inv_4 Z_4 out_4 vdd gnd pinv_6
Xpre_nand_inv_5 Z_5 out_5 vdd gnd pinv_6
Xpre_nand_inv_6 Z_6 out_6 vdd gnd pinv_6
Xpre_nand_inv_7 Z_7 out_7 vdd gnd pinv_6
XXpre3x8_nand_0 inbar_0 inbar_1 inbar_2 Z_0 vdd gnd pnand3_1
XXpre3x8_nand_1 in_0 inbar_1 inbar_2 Z_1 vdd gnd pnand3_1
XXpre3x8_nand_2 inbar_0 in_1 inbar_2 Z_2 vdd gnd pnand3_1
XXpre3x8_nand_3 in_0 in_1 inbar_2 Z_3 vdd gnd pnand3_1
XXpre3x8_nand_4 inbar_0 inbar_1 in_2 Z_4 vdd gnd pnand3_1
XXpre3x8_nand_5 in_0 inbar_1 in_2 Z_5 vdd gnd pnand3_1
XXpre3x8_nand_6 inbar_0 in_1 in_2 Z_6 vdd gnd pnand3_1
XXpre3x8_nand_7 in_0 in_1 in_2 Z_7 vdd gnd pnand3_1
.ENDS hierarchical_predecode3x8_1

.SUBCKT bank dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 rbl_bl_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 addr0_9 s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: dout0_8 
* OUTPUT: dout0_9 
* OUTPUT: dout0_10 
* OUTPUT: dout0_11 
* OUTPUT: dout0_12 
* OUTPUT: dout0_13 
* OUTPUT: dout0_14 
* OUTPUT: dout0_15 
* OUTPUT: dout0_16 
* OUTPUT: dout0_17 
* OUTPUT: dout0_18 
* OUTPUT: dout0_19 
* OUTPUT: dout0_20 
* OUTPUT: dout0_21 
* OUTPUT: dout0_22 
* OUTPUT: dout0_23 
* OUTPUT: dout0_24 
* OUTPUT: dout0_25 
* OUTPUT: dout0_26 
* OUTPUT: dout0_27 
* OUTPUT: dout0_28 
* OUTPUT: dout0_29 
* OUTPUT: dout0_30 
* OUTPUT: dout0_31 
* OUTPUT: rbl_bl_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : din0_8 
* INPUT : din0_9 
* INPUT : din0_10 
* INPUT : din0_11 
* INPUT : din0_12 
* INPUT : din0_13 
* INPUT : din0_14 
* INPUT : din0_15 
* INPUT : din0_16 
* INPUT : din0_17 
* INPUT : din0_18 
* INPUT : din0_19 
* INPUT : din0_20 
* INPUT : din0_21 
* INPUT : din0_22 
* INPUT : din0_23 
* INPUT : din0_24 
* INPUT : din0_25 
* INPUT : din0_26 
* INPUT : din0_27 
* INPUT : din0_28 
* INPUT : din0_29 
* INPUT : din0_30 
* INPUT : din0_31 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : addr0_8 
* INPUT : addr0_9 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xreplica_bitcell_array bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 rbl_bl_0 rbl_br_0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 wl_en0 vdd gnd replica_bitcell_array_0
Xport_data0 rbl_bl_0 rbl_br_0 bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62 br_62 bl_63 br_63 bl_64 br_64 bl_65 br_65 bl_66 br_66 bl_67 br_67 bl_68 br_68 bl_69 br_69 bl_70 br_70 bl_71 br_71 bl_72 br_72 bl_73 br_73 bl_74 br_74 bl_75 br_75 bl_76 br_76 bl_77 br_77 bl_78 br_78 bl_79 br_79 bl_80 br_80 bl_81 br_81 bl_82 br_82 bl_83 br_83 bl_84 br_84 bl_85 br_85 bl_86 br_86 bl_87 br_87 bl_88 br_88 bl_89 br_89 bl_90 br_90 bl_91 br_91 bl_92 br_92 bl_93 br_93 bl_94 br_94 bl_95 br_95 bl_96 br_96 bl_97 br_97 bl_98 br_98 bl_99 br_99 bl_100 br_100 bl_101 br_101 bl_102 br_102 bl_103 br_103 bl_104 br_104 bl_105 br_105 bl_106 br_106 bl_107 br_107 bl_108 br_108 bl_109 br_109 bl_110 br_110 bl_111 br_111 bl_112 br_112 bl_113 br_113 bl_114 br_114 bl_115 br_115 bl_116 br_116 bl_117 br_117 bl_118 br_118 bl_119 br_119 bl_120 br_120 bl_121 br_121 bl_122 br_122 bl_123 br_123 bl_124 br_124 bl_125 br_125 bl_126 br_126 bl_127 br_127 bl_128 br_128 bl_129 br_129 bl_130 br_130 bl_131 br_131 bl_132 br_132 bl_133 br_133 bl_134 br_134 bl_135 br_135 bl_136 br_136 bl_137 br_137 bl_138 br_138 bl_139 br_139 bl_140 br_140 bl_141 br_141 bl_142 br_142 bl_143 br_143 bl_144 br_144 bl_145 br_145 bl_146 br_146 bl_147 br_147 bl_148 br_148 bl_149 br_149 bl_150 br_150 bl_151 br_151 bl_152 br_152 bl_153 br_153 bl_154 br_154 bl_155 br_155 bl_156 br_156 bl_157 br_157 bl_158 br_158 bl_159 br_159 bl_160 br_160 bl_161 br_161 bl_162 br_162 bl_163 br_163 bl_164 br_164 bl_165 br_165 bl_166 br_166 bl_167 br_167 bl_168 br_168 bl_169 br_169 bl_170 br_170 bl_171 br_171 bl_172 br_172 bl_173 br_173 bl_174 br_174 bl_175 br_175 bl_176 br_176 bl_177 br_177 bl_178 br_178 bl_179 br_179 bl_180 br_180 bl_181 br_181 bl_182 br_182 bl_183 br_183 bl_184 br_184 bl_185 br_185 bl_186 br_186 bl_187 br_187 bl_188 br_188 bl_189 br_189 bl_190 br_190 bl_191 br_191 bl_192 br_192 bl_193 br_193 bl_194 br_194 bl_195 br_195 bl_196 br_196 bl_197 br_197 bl_198 br_198 bl_199 br_199 bl_200 br_200 bl_201 br_201 bl_202 br_202 bl_203 br_203 bl_204 br_204 bl_205 br_205 bl_206 br_206 bl_207 br_207 bl_208 br_208 bl_209 br_209 bl_210 br_210 bl_211 br_211 bl_212 br_212 bl_213 br_213 bl_214 br_214 bl_215 br_215 bl_216 br_216 bl_217 br_217 bl_218 br_218 bl_219 br_219 bl_220 br_220 bl_221 br_221 bl_222 br_222 bl_223 br_223 bl_224 br_224 bl_225 br_225 bl_226 br_226 bl_227 br_227 bl_228 br_228 bl_229 br_229 bl_230 br_230 bl_231 br_231 bl_232 br_232 bl_233 br_233 bl_234 br_234 bl_235 br_235 bl_236 br_236 bl_237 br_237 bl_238 br_238 bl_239 br_239 bl_240 br_240 bl_241 br_241 bl_242 br_242 bl_243 br_243 bl_244 br_244 bl_245 br_245 bl_246 br_246 bl_247 br_247 bl_248 br_248 bl_249 br_249 bl_250 br_250 bl_251 br_251 bl_252 br_252 bl_253 br_253 bl_254 br_254 bl_255 br_255 dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 dout0_8 dout0_9 dout0_10 dout0_11 dout0_12 dout0_13 dout0_14 dout0_15 dout0_16 dout0_17 dout0_18 dout0_19 dout0_20 dout0_21 dout0_22 dout0_23 dout0_24 dout0_25 dout0_26 dout0_27 dout0_28 dout0_29 dout0_30 dout0_31 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7 din0_8 din0_9 din0_10 din0_11 din0_12 din0_13 din0_14 din0_15 din0_16 din0_17 din0_18 din0_19 din0_20 din0_21 din0_22 din0_23 din0_24 din0_25 din0_26 din0_27 din0_28 din0_29 din0_30 din0_31 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4 sel0_5 sel0_6 sel0_7 s_en0 p_en_bar0 w_en0 vdd gnd port_data_0
Xport_address0 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 addr0_8 addr0_9 wl_en0 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 wl_89 wl_90 wl_91 wl_92 wl_93 wl_94 wl_95 wl_96 wl_97 wl_98 wl_99 wl_100 wl_101 wl_102 wl_103 wl_104 wl_105 wl_106 wl_107 wl_108 wl_109 wl_110 wl_111 wl_112 wl_113 wl_114 wl_115 wl_116 wl_117 wl_118 wl_119 wl_120 wl_121 wl_122 wl_123 wl_124 wl_125 wl_126 wl_127 vdd gnd port_address_0
Xcol_address_decoder0 addr0_0 addr0_1 addr0_2 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4 sel0_5 sel0_6 sel0_7 vdd gnd hierarchical_predecode3x8_1
.ENDS bank

* ptx M{0} {1} pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_7 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_7

* ptx M{0} {1} nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p

* ptx M{0} {1} pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p

.SUBCKT pinv_8 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.54u l=0.05u pd=1.18u ps=1.18u as=0.07p ad=0.07p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pinv_8

.SUBCKT dff_buf_0 D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff D qint clk vdd gnd dff
Xdff_buf_inv1 qint Qb vdd gnd pinv_7
Xdff_buf_inv2 Qb Q vdd gnd pinv_8
.ENDS dff_buf_0

.SUBCKT dff_buf_array_0 din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_r0_c0 din_0 dout_0 dout_bar_0 clk vdd gnd dff_buf_0
Xdff_r1_c0 din_1 dout_1 dout_bar_1 clk vdd gnd dff_buf_0
.ENDS dff_buf_array_0

.SUBCKT pnand2_1 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.02p ad=0.02p
.ENDS pnand2_1

.SUBCKT pinv_9 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_9

.SUBCKT pdriver_1 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 4]
Xbuf_inv1 A Zb1_int vdd gnd pinv_9
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_9
Xbuf_inv3 Zb2_int Z vdd gnd pinv_8
.ENDS pdriver_1

.SUBCKT pand2_0 A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand2_nand A B zb_int vdd gnd pnand2_1
Xpand2_inv zb_int Z vdd gnd pdriver_1
.ENDS pand2_0

* ptx M{0} {1} nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p

.SUBCKT pinv_10 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=21 w=0.8225u l=0.05u pd=1.75u ps=1.75u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=21 w=0.275u l=0.05u pd=0.65u ps=0.65u as=0.03p ad=0.03p
.ENDS pinv_10

* ptx M{0} {1} nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p

.SUBCKT pinv_11 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=81 w=0.8525u l=0.05u pd=1.81u ps=1.81u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=81 w=0.28500000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_11

.SUBCKT pbuf_0 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1 A zb_int vdd gnd pinv_10
Xbuf_inv2 zb_int Z vdd gnd pinv_11
.ENDS pbuf_0

* ptx M{0} {1} nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_12 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_12

* ptx M{0} {1} nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_13 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_13

* ptx M{0} {1} nmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=9 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p

.SUBCKT pinv_14 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.81u l=0.05u pd=1.72u ps=1.72u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
.ENDS pinv_14

* ptx M{0} {1} nmos_vtg m=26 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=26 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p

.SUBCKT pinv_15 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=26 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=26 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p
.ENDS pinv_15

.SUBCKT pdriver_2 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 27, 80]
Xbuf_inv1 A Zb1_int vdd gnd pinv_9
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_9
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_12
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_13
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_14
Xbuf_inv6 Zb5_int Z vdd gnd pinv_15
.ENDS pdriver_2

* ptx M{0} {1} nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p

.SUBCKT pinv_16 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.675u l=0.05u pd=1.45u ps=1.45u as=0.08p ad=0.08p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.225u l=0.05u pd=0.55u ps=0.55u as=0.03p ad=0.03p
.ENDS pinv_16

* ptx M{0} {1} nmos_vtg m=5 w=0.2525u l=0.05u pd=0.60u ps=0.60u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=5 w=0.755u l=0.05u pd=1.61u ps=1.61u as=0.09p ad=0.09p

.SUBCKT pinv_17 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=5 w=0.755u l=0.05u pd=1.61u ps=1.61u as=0.09p ad=0.09p
Mpinv_nmos Z A gnd gnd nmos_vtg m=5 w=0.2525u l=0.05u pd=0.60u ps=0.60u as=0.03p ad=0.03p
.ENDS pinv_17

* ptx M{0} {1} nmos_vtg m=14 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=14 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p

.SUBCKT pinv_18 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=14 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=14 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p
.ENDS pinv_18

.SUBCKT pdriver_3 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 2, 5, 14, 43]
Xbuf_inv1 A Zb1_int vdd gnd pinv_9
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_9
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_7
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_16
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_17
Xbuf_inv6 Zb5_int Z vdd gnd pinv_18
.ENDS pdriver_3

* ptx M{0} {1} nmos_vtg m=13 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=13 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p

.SUBCKT pinv_19 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=13 w=0.8300000000000001u l=0.05u pd=1.76u ps=1.76u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=13 w=0.2775u l=0.05u pd=0.66u ps=0.66u as=0.03p ad=0.03p
.ENDS pinv_19

.SUBCKT pand3_0 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_19
.ENDS pand3_0

* ptx M{0} {1} nmos_vtg m=11 w=0.2625u l=0.05u pd=0.62u ps=0.62u as=0.03p ad=0.03p

* ptx M{0} {1} pmos_vtg m=11 w=0.785u l=0.05u pd=1.67u ps=1.67u as=0.10p ad=0.10p

.SUBCKT pinv_20 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=11 w=0.785u l=0.05u pd=1.67u ps=1.67u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=11 w=0.2625u l=0.05u pd=0.62u ps=0.62u as=0.03p ad=0.03p
.ENDS pinv_20

.SUBCKT pand3_1 A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpand3_nand A B C zb_int vdd gnd pnand3_1
Xpand3_inv zb_int Z vdd gnd pinv_20
.ENDS pand3_1

* ptx M{0} {1} nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p

.SUBCKT pinv_21 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=9 w=0.84u l=0.05u pd=1.78u ps=1.78u as=0.10p ad=0.10p
Mpinv_nmos Z A gnd gnd nmos_vtg m=9 w=0.28u l=0.05u pd=0.66u ps=0.66u as=0.04p ad=0.04p
.ENDS pinv_21

* ptx M{0} {1} nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p

* ptx M{0} {1} pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p

.SUBCKT pinv_22 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=27 w=0.85u l=0.05u pd=1.80u ps=1.80u as=0.11p ad=0.11p
Mpinv_nmos Z A gnd gnd nmos_vtg m=27 w=0.28250000000000003u l=0.05u pd=0.67u ps=0.67u as=0.04p ad=0.04p
.ENDS pinv_22

.SUBCKT pdriver_4 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 3, 9, 28, 85]
Xbuf_inv1 A Zb1_int vdd gnd pinv_9
Xbuf_inv2 Zb1_int Zb2_int vdd gnd pinv_9
Xbuf_inv3 Zb2_int Zb3_int vdd gnd pinv_12
Xbuf_inv4 Zb3_int Zb4_int vdd gnd pinv_13
Xbuf_inv5 Zb4_int Zb5_int vdd gnd pinv_21
Xbuf_inv6 Zb5_int Z vdd gnd pinv_22
.ENDS pdriver_4

.SUBCKT pinv_23 A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03p ad=0.03p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01p ad=0.01p
.ENDS pinv_23

.SUBCKT delay_chain_0 in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0 in dout_1 vdd gnd pinv_23
Xdload_0_0 dout_1 n_0_0 vdd gnd pinv_23
Xdload_0_1 dout_1 n_0_1 vdd gnd pinv_23
Xdload_0_2 dout_1 n_0_2 vdd gnd pinv_23
Xdload_0_3 dout_1 n_0_3 vdd gnd pinv_23
Xdinv1 dout_1 dout_2 vdd gnd pinv_23
Xdload_1_0 dout_2 n_1_0 vdd gnd pinv_23
Xdload_1_1 dout_2 n_1_1 vdd gnd pinv_23
Xdload_1_2 dout_2 n_1_2 vdd gnd pinv_23
Xdload_1_3 dout_2 n_1_3 vdd gnd pinv_23
Xdinv2 dout_2 dout_3 vdd gnd pinv_23
Xdload_2_0 dout_3 n_2_0 vdd gnd pinv_23
Xdload_2_1 dout_3 n_2_1 vdd gnd pinv_23
Xdload_2_2 dout_3 n_2_2 vdd gnd pinv_23
Xdload_2_3 dout_3 n_2_3 vdd gnd pinv_23
Xdinv3 dout_3 dout_4 vdd gnd pinv_23
Xdload_3_0 dout_4 n_3_0 vdd gnd pinv_23
Xdload_3_1 dout_4 n_3_1 vdd gnd pinv_23
Xdload_3_2 dout_4 n_3_2 vdd gnd pinv_23
Xdload_3_3 dout_4 n_3_3 vdd gnd pinv_23
Xdinv4 dout_4 dout_5 vdd gnd pinv_23
Xdload_4_0 dout_5 n_4_0 vdd gnd pinv_23
Xdload_4_1 dout_5 n_4_1 vdd gnd pinv_23
Xdload_4_2 dout_5 n_4_2 vdd gnd pinv_23
Xdload_4_3 dout_5 n_4_3 vdd gnd pinv_23
Xdinv5 dout_5 dout_6 vdd gnd pinv_23
Xdload_5_0 dout_6 n_5_0 vdd gnd pinv_23
Xdload_5_1 dout_6 n_5_1 vdd gnd pinv_23
Xdload_5_2 dout_6 n_5_2 vdd gnd pinv_23
Xdload_5_3 dout_6 n_5_3 vdd gnd pinv_23
Xdinv6 dout_6 dout_7 vdd gnd pinv_23
Xdload_6_0 dout_7 n_6_0 vdd gnd pinv_23
Xdload_6_1 dout_7 n_6_1 vdd gnd pinv_23
Xdload_6_2 dout_7 n_6_2 vdd gnd pinv_23
Xdload_6_3 dout_7 n_6_3 vdd gnd pinv_23
Xdinv7 dout_7 dout_8 vdd gnd pinv_23
Xdload_7_0 dout_8 n_7_0 vdd gnd pinv_23
Xdload_7_1 dout_8 n_7_1 vdd gnd pinv_23
Xdload_7_2 dout_8 n_7_2 vdd gnd pinv_23
Xdload_7_3 dout_8 n_7_3 vdd gnd pinv_23
Xdinv8 dout_8 out vdd gnd pinv_23
Xdload_8_0 out n_8_0 vdd gnd pinv_23
Xdload_8_1 out n_8_1 vdd gnd pinv_23
Xdload_8_2 out n_8_2 vdd gnd pinv_23
Xdload_8_3 out n_8_3 vdd gnd pinv_23
.ENDS delay_chain_0

.SUBCKT control_logic_rw csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* word_size 32
Xctrl_dffs csb web cs_bar cs we_bar we clk_buf vdd gnd dff_buf_array_0
Xclkbuf clk clk_buf vdd gnd pdriver_2
Xinv_clk_bar clk_buf clk_bar vdd gnd pinv_9
Xand2_gated_clk_bar cs clk_bar gated_clk_bar vdd gnd pand2_0
Xand2_gated_clk_buf clk_buf cs gated_clk_buf vdd gnd pand2_0
Xbuf_wl_en gated_clk_bar wl_en vdd gnd pdriver_3
Xrbl_bl_delay_inv rbl_bl_delay rbl_bl_delay_bar vdd gnd pinv_9
Xw_en_and we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd pand3_0
Xbuf_s_en_and rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd pand3_1
Xdelay_chain rbl_bl rbl_bl_delay vdd gnd delay_chain_0
Xnand_p_en_bar gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd pnand2_1
Xbuf_p_en_bar p_en_bar_unbuf p_en_bar vdd gnd pdriver_4
.ENDS control_logic_rw

.SUBCKT sram_32_1024_freepdk45 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] csb0 web0 clk0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : din0[8] 
* INPUT : din0[9] 
* INPUT : din0[10] 
* INPUT : din0[11] 
* INPUT : din0[12] 
* INPUT : din0[13] 
* INPUT : din0[14] 
* INPUT : din0[15] 
* INPUT : din0[16] 
* INPUT : din0[17] 
* INPUT : din0[18] 
* INPUT : din0[19] 
* INPUT : din0[20] 
* INPUT : din0[21] 
* INPUT : din0[22] 
* INPUT : din0[23] 
* INPUT : din0[24] 
* INPUT : din0[25] 
* INPUT : din0[26] 
* INPUT : din0[27] 
* INPUT : din0[28] 
* INPUT : din0[29] 
* INPUT : din0[30] 
* INPUT : din0[31] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : addr0[8] 
* INPUT : addr0[9] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* OUTPUT: dout0[8] 
* OUTPUT: dout0[9] 
* OUTPUT: dout0[10] 
* OUTPUT: dout0[11] 
* OUTPUT: dout0[12] 
* OUTPUT: dout0[13] 
* OUTPUT: dout0[14] 
* OUTPUT: dout0[15] 
* OUTPUT: dout0[16] 
* OUTPUT: dout0[17] 
* OUTPUT: dout0[18] 
* OUTPUT: dout0[19] 
* OUTPUT: dout0[20] 
* OUTPUT: dout0[21] 
* OUTPUT: dout0[22] 
* OUTPUT: dout0[23] 
* OUTPUT: dout0[24] 
* OUTPUT: dout0[25] 
* OUTPUT: dout0[26] 
* OUTPUT: dout0[27] 
* OUTPUT: dout0[28] 
* OUTPUT: dout0[29] 
* OUTPUT: dout0[30] 
* OUTPUT: dout0[31] 
* POWER : vdd 
* GROUND: gnd 
Xbank0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30] dout0[31] rbl_bl0 bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] a0[0] a0[1] a0[2] a0[3] a0[4] a0[5] a0[6] a0[7] a0[8] a0[9] s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd bank
Xcontrol0 csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd control_logic_rw
Xrow_address0 addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr0[8] addr0[9] a0[3] a0[4] a0[5] a0[6] a0[7] a0[8] a0[9] clk_buf0 vdd gnd row_addr_dff
Xcol_address0 addr0[0] addr0[1] addr0[2] a0[0] a0[1] a0[2] clk_buf0 vdd gnd col_addr_dff
Xdata_dff0 din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23] din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] bank_din0[0] bank_din0[1] bank_din0[2] bank_din0[3] bank_din0[4] bank_din0[5] bank_din0[6] bank_din0[7] bank_din0[8] bank_din0[9] bank_din0[10] bank_din0[11] bank_din0[12] bank_din0[13] bank_din0[14] bank_din0[15] bank_din0[16] bank_din0[17] bank_din0[18] bank_din0[19] bank_din0[20] bank_din0[21] bank_din0[22] bank_din0[23] bank_din0[24] bank_din0[25] bank_din0[26] bank_din0[27] bank_din0[28] bank_din0[29] bank_din0[30] bank_din0[31] clk_buf0 vdd gnd data_dff
.ENDS sram_32_1024_freepdk45
