`include "../common/packet_in.sv"
`include "../common/packet_out.sv"
`include "../add/sequence_in.sv"
`include "../add/fsm_add.sv"
`include "../common/sequencer.sv"
`include "../common/driver.sv"
`include "../common/driver_out.sv"
`include "../common/monitor.sv"
`include "../common/monitor_out.sv"
`include "../common/agent.sv"
`include "../common/agent_out.sv"
`include "../add/refmod.sv"
`include "../common/comparator.sv"
`include "../common/env.sv"
`include "../common/simple_test.sv"
`include "../src/adder.sv"